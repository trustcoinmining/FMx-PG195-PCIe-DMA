`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
eXm8mGGNxF6S7JgSE9KR4pzbZ3WeLCvd1Qpi4ZqeT3EcGZgcTjif8pyb/o3+ZI6R3oU6rEMUYPFu
qEa8XwfdfQ==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
S9DWlcj0qvlNCDKyR5+ELekKiEo44BcOStsDOJx0v2NVuGcg2+04VEW1g1HWZMCh4OxUq61m78q1
0Kn0CqzIZu2qHvUoU93VN9i7zrXOwMNK9MyWDRE65jMgRzDDXsFfL3G8/jDxiCGn9OHJF+T06GJR
X8TLmy5iQdI67oP5Eq8=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y5dHosYSgCHMyWKz7ujToKtCGB0s1lJTDuynh01WO11DzbFG8RPWUBMp7XLEfr4hCYhNkQ7m3jJk
VUgle22Kh7D0/kGhoarCi6ym9oqRQHT7PXQmIEqu63vLrFam70rxUTGkShMESadKCm0cElHJjRJT
hlCvgwcm/4uim6dJGmQvf9h8auBnUmRrV9ibmkjC9Y+BFvMR/BPr4d32opmVnV/Yy9TEIf2j3nml
pSRZkWiZwR9KiYVy+9nLju154KCezlqCOUIDT2kcE55OFk+e1fj7d740rgviVDbCi2uTCd4sm7Gd
wVjR1yIA9oXSArcXfN+nPxzpC/itZLYqXuV6Eg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QQduTFGip3mKvMV++cB5PQonf7i+fhZYzaWPONWWgXaFzn3WW4r9gb+BwTGuqZjKe7kkfaA8e2H3
rI1IgppKW9MGHRZ+Gvjenf0m9y7tFVQXmclPgb6iI4E5MH54XJYsx9pFPLcGosui6Mo8C7iKcSnL
GCmvskWnuO+IGcshduWu1PVn/Oz+E6dSRaOmHnIMvun/rQ/Bi7mBHaB1/YQRB8ND8zWM1TmfsWgI
2d7LjLnZMPoqQuTpECzal7DxSCXSWI+17PZOOHzwiz5QGoHDLKO/+fzGIgV10IBhczOYtwJIOTk1
AQnv02ybkp2SCMKq2d2UpMezuUgNN3Qi6+iFdg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W+V3hT9NuKxb/1LWlhZ8Tixa3j0ef5yysCyYpdj4Bpe9o5XW3AlaBsVBMW5aoTShMTHI4m5kUD3k
ojMb6Le0vKYs1TV0AMrgmD+oGSwajLcWvcfmJy10GPagtygmNDl7DDJkHrVquJpRjOvGqNvdWugO
gTZhB5gmTXbT8RXvr1jnb5q5/qHBYpiFyojNOM+0wr4tcbZyzbmcWVgdKdPs9AtOeXrFChoBNKzO
ZfDiVshP70IL+hqQownr9okwDrx/bq0eRyJF8lJivvIyNKC1HOu4C9kIvFcPv/sEqvYuCFolRkSn
OP5fjmiQAdrkkd73H05nJlVhgar08HIq4tiX8Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ipNpLEzwh2bJzRySQ+x8H8oCxhmvdEl5+u9ySbaCMJQlxTPTA20LakbPY6DFOu+SXAVpf7hsqqa6
rNoFKs3gmpQdD438VCVjCE5egTKa6GOihOwoe6eUDBJ6QU3cnpjYIHgycGnbwjcD22PBThvQ+SNR
RL9xggQu3H51RiP/vHo=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RuOz8zdtGw7N501KzSeNo1+Gl58MGQrvQybU+QuHBPIm/+ZQwjx1xd6wL4ZfwhWrX0YXB3JBdVLx
3qCtjufI5dyfBmIUGRctH0JuJEE5EtjvN1dS4sUcx1JQpqw32E+RMCPNy2LWSRjLi+gfXOSiv2tk
RbQA4lXoJPY7YnFsLPBn91jSdoHpZo2A9m/oCXgI5IObyf/3ytESVvI9kMIj2yVpvun48/zGB6NO
sMrk54Q2bUTuNA1Ylc53OU2gRT0MGNb//mrPxPAVewZWBY1z74+Y5fBKKB4q6ZidjkvokF/1UYz0
97VTxNPtC59z/+8+Deqo/osa57sAFVXmVegb2g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1051216)
`protect data_block
Oy6MSkudSG0mKc+cpvU3rRghbLKhjAz/Oe1ZR5uU4al24QXNJESLqPiy6RlzaVvgqD4yU+9h9PlZ
7xtnz5sbynohOVsiE7BpyMQyZsmDxGtuML2v/eKpxoct465329cOTJpT2nNFotqmyDZzU4ajthC9
RUY6h+TW7VuP4EBbcVb/hZHPngrl44nvY1XcJL48G0Xw0gMCnOrktsqjAZwGLlK/533SY1ftgPOZ
bn6wc1QrzuAe5PJLrMxHB/e2K8W58hbk0eucjT9kUKUfq1OrOGm63N2FeFxxtNG7CfGBOtSWWt2O
B49b3R9GlXm2YmgiK+VA7u6rI53/6USry/nTyQIo9b8EW+4jBn7+reU175Lo2yEUReBlhk8sDN3q
mBKHy7n/c7wNX9KhdsUofokZt9JcINXJ7ZnI/o35PZEqs5dYMNzF2qlGQfYUtLnhyGJlR0Leztbs
BlJkxTqboNH/+VJ6gYEAIRWm93ARkn/ZQJFiTRS4eyhQFm40j0eI4D0jOqlokTy6pYe8ts1g1B2o
2fBrWZYoO9d1xIwLyqaxTa9ol1C2+qUrprP9EkTTWH4Ejqa3qnZy5TT0YE58Gc6E2T8/0qbJkMBc
JpMlk8l4Lb/US2aSaZ374RqFVHnnLojOTMvf1aZf8bze/VI2LpO64Life0W2HINgDSOrx2dfs7WX
5//Jd6z5AjHvaSIEryTblDQZT3u4UC7tSYlAksdmyZRU62ZgtLhVhrj8GFMnkyMt5L/VrMChdzVd
yi4QJ7gUHOKtBOk5bY5iJkmDfJKLbvyfPT869QkucxJK1v57NUnnmVYP245sneJEd+2mbtzO8vDl
5PQDbmtjDcbOQYScCdOPnzZvK90XMzjm7+bgJhENkEePg2idZCnhJIpl5z4St1YdmUHMacraGsF5
AvcG4EylEDL3YwZFT3c65CmL7k5iSDD7ItYsMvKVQ6kgHS2Km4jJr4+vGOUkxMRMDgxjouQwsPBc
MYPtUCo5r54DhyOnozpupN2jzkOiK9bPEnKHkHIXLVUdpjST8VN1j8y1+E1Lydt7ycP1UoomKWym
G0YwbyVX0J7w/gDKYJ/+edhR4p3LYXIEAwRz4ljpoEwTqhfprUwTG+2w6TJeE2Kn02bRTkwR6YC8
yM0CY3JZG0BZ56uJ7ogm2GsRv7F062pOfXPhv5BF+9M0Xlr5Uk9JaV3ngoGOo0Fih13huH+27kro
hc1AuT404DFCbXkIwEdKejs3y7v5ZUeo01beh/pJlCPpk/8bjBMVhKWeDOvbJ2jv0wTYC2SGAwx3
FqLwuOECcNsgW8Zx7iJEgSWTgj4UiJboXSTB1fc17T8SMJ0F8DqoI3KcMwSgas2fRE3qDWr8Pi7v
tIK+GcnmbneV8tSCxoCJDlMK6y6ij1VUSGbCPLfBEZ23M7qRzN06SbP7eaxH8dA2jGbk9vjO05jg
m7/IYEHs94jLat1qQwzLCT961lbP4a1yyW1NewFWQ+7g4++Kwvr2wapYVsHlhz9RF0jNDQ8EEXqF
Y+C97t/OZUCNiountEJQaOel9K/SK2Rcfx80SSnorzF6f8jtBSaGezXUBM+TnuPRoZBwY5YgZZIr
Bttzli0AbeCcmEe5ECF9LikWKZOgouAzfGN8fMliFsaOsKZ4lD9fyU4NcDhZRaqT+vwpWOYrmW33
7rVIYjmHPgtw48UkI9ZRWb3WfM74/iSpAT5Wm8EiF+FWQtXFplspQWdOTqyZ39zFCwxjX5M+qx4+
l1nkUQLCIzGWV6AfaVZpzsCnc8AMqfIBHPx9qW9PcTI2oF2cUe/DoC3olIwCrfOc1m2TMTkqbxOO
q1BBqGVSwX5WnSiuplhFRAox/HM1FdKLranpXAuQpBDvTfNjmVi1rTOP3I5+RIOHUIHHYR3TU1SZ
ThXcoSMcGDeDNHSjFN1oI87pD4nZpchlGCHusSC2QDp9KiXIybYtb6SUZh8CPxSrEfcLgfhA4gCE
s5fKtBJdh0Wb+kEXoQhUBDnXg+4QA4kJWAVPImCkeCFYqF42jIDauhjjf8qNhI5avmmh4wS02H6j
JgkQ218AmIos0XpgmAcyoo/iLAPYaOmL6XInpa/u10KqwQJ5wOHzZd8XD+Zq+q3RlTbwZ9sJpmZX
S3cxVE/pHTlHWfx5wp4ZmLrnmjuXzGNBd2Mf8R6uS90no8XPgj2MDuCiD5XKg97FD7xXDAt6yPBR
1VdoDWc2VZZEaVe7wpwffSTXY54/S9hTxJROH5ttCCM2ZU9EIDuo4J0CVBTUiIy+v629m10BYGFk
BD85UEGOJXei+nOniGOfeY/nYfreqwrQEeeWe3cRmAs62A3uk3N+FhXv9kAVKPD9kRbxla2uBGBB
UoUSBF6U1qKw1zSabz205u6bPcfPwQ0mpbFXpkxjnqPZ40YqbZ9NInU6LpuroJptxhcT6M/2i+fW
s6UNsqHWrLbPZ1DcRaLxntfWfiagSvrgtcR9jqjoStO9SFHDAf+CsvvNKHmBKXEsoZR1PATIpLl1
4qDKQUNGJCxwAOLgv82mPuZHVywMgtBrvJALx3ODmtemYcQlE8rMaSsObHqVZ/Tyr/m8y77yY59K
YxyvAzTLFZ2Vkp7Sleh2hWGjxQWv9Nm1zDKfyE2vubApsI1qCKkvX+MZ/C4pTRAKyAk42FJi5Yan
xhmEWamjddrW0x/3pV7serzb4M9Yw6rEjDYZFobDs2e6VxmYQOLVIJMQe8DWXEcRU/66e4aYp0Zd
OTIPQdYcva8uSnxvw1OeIEOUhnOmcfalgNTJOejMQOKzfg6ljCZ1P3cKAmqxwWjzlcaxyrtaVbBO
0p9xQG8xeK1IgS21FbMAFEcIBlTJcnHaES4tBbfgjyRt2x5A+9MLLtZClOuvyGbkB4F48MP4/w+W
g7XLZejlPQmCV/GLyJnnWdlFJeoi3m5vo3GPbOddeisSwzLPEwDbMmWD7OrTDMz0KNP/gsGIWeYP
j5i18GK+uCYOgCuqymmy6UmvYwNSXMUlfxzGtgRxTuoEIrCcxAvLargCe8hNJTqMZUrmgs9fRcZ1
OQv/dExFVVXj62MZ7cOVQwT6cJQBdAT/zq9V5pmPo2JjiZ3pHqN8aZB19SqQGhhPehgcDZAg97CO
6CmBz2ddDmjPwOo4IU1ikOM0er0AOzs7vW7A3whKDPH9V3ZBYxCVO6FKS9dLG4qwkkMUftl9ursn
ZvWrrsAdwUr8BpTItLjzEMBKkkswMSJWAlVpYCVdKIFttPaA9pSV1kTHnnnpJD4mkULGU71q5nD0
TaDXfVc5raVauxJffNWzg/vEYuv01uOYjmeCsRH/X2Y3wwb/SWe+Nwds3ZcALn1+WF4aDA4xs1/v
tVa7K3GuEy5O2iAwOwFLxErDl91Vx4cSLf+XvuhXY11v8VHUrkTGYBOlxgoB7LHUMx2wYFff5CDX
Nf+h7PRXnp4/dCEOSPk4EjaVY5yjgGRjF2nQIZ1O6EJA+zmDi7U9nqJkAVBLgeWsRQJXth/XPBmT
6+HRcej58RqTZymBEVltZTtqD4B1KZJAgzDOsy1wWu+aZRaZ0qkZk/4ITyXHVxSqdfQsjAiJgTxU
byMfUHsTjK3WouSiDKm268OrgpYqMXaki3cTQPJK9YJGayhBBz9lFEX/fgC2LnGKTJ/w+C05njBA
QNiRlJYdZ5madRyc72QQWP1JffBoKGDxUCgFJXga+vJJvIPEnRjk3fxC9x8+/7uoINOX88k/dcc5
E0I48a0SKJBmEBHmLt93Hq7IyWCvKQgDMSBAGpUtF6TSCGLJxf8KnvEVwcRN64F+xxvDcJZJ+y4C
d8+GVY+MkKIJGf8j3DGE6cXIbvWPRBXBhDCGTRk7BdDviXphxPuCPZqwEhfht5SYHnRrZkKrPGp5
ti+091OQ7ez8ArQYhjHcrYrqBfYcWSlvahlIv2brb+Y97BEgKGZBCa4nNFDXVulG6iPRjwvVVIQZ
JrmYGcPtGSgYJPylnoRq0kwUPcVsSrCr2WvJwRRcayxDJ0tKk1IIe2SqVqZYyk+5SpxdSH9dhjsO
3hz6wWpsxFGfxE3ErU1XTnw8TIqQ9EUTWv7lsF4Qj6yDRz2FoBn1+xeicQzvGob9skCspXEXL/pg
fNHeQruQW+9xO8qUUWzI1GurNmop7qIRq3djNJDfdtJ7m0Mmav1wU+8A2qUaLTse8lX1nxTqAuZ3
0cwB1whvLVdJ062sDb43rXrmMxpgxltvS3/Lm4HUsV66qZDoLq86g+41lkCTa9ignWWqkatqPjRb
koWDUis4zCyg5rRUxGOOw3s7u1bHhiyvv2sJ8dgeKOulQ7Rs+kixZ9EHoBJgOm7kiEvwJO4REmy9
gq3vcZiwi17TtJ2XpEd4D/Run1nMPRmpkZDm2FwfRGwYTwlhDdV7towCK3EgpxcGAxIQ46gVxtU/
Iy3x41w4KP7dkUKpe2lekJ5ldgj7FdmHPyYP+pN2YmOYUP6gbKTtrhvw/4obfHELx9DbrTMJppzK
3qGMZsrddkduADLBaI/4VQZKtDZLO0eKCCdOU/z6u/F+Q+FxsO2gjF6iAb9Gs795lsFTC4/nPd5G
MngCl3IsavsRBxwXigSAlvq68cJzBLb+AE6SEOsFXSzy0Tm3kf12Xf08VrT9IEVafq9j0R3fXagE
s+6XF6TB7C67le2g8GjkxPgfF3N3dJLmgoSVlAqBPvsgRhmXn4Tm+Ij6dYPscz7sruyVhh6TRnfS
IuRq8S2OSf/CcNw2uyhOs4UF6gEA9uV4x8MZ63XtNyMzQloU3jsq5jwZc/HmLQmd5K478xCVgiIe
NgPNsfMDvFFLLxJBIcR7RVRHXImKpNLROF05efnrwFAeGrcuA6I4bnzJjoaimJyG/ke+WYDxmdn+
VrFrYy4ezYak7FY4xZZChiQ/MTyNw7/BlejklEHZzyfNvdJMgPlxa75pXNZKYS0kCQRjvOipVCN5
/hilmnespLg1ofb2voBMH5/8f6+924sud7IV6YEgt4+FSQs1ZxwUgPXa0SXMuf8L55hjYbkyIUhc
BsXaRBeQFDFLxtRusJ7NuJLuDy8tbn8CwZxgqqA7W5qFes9LMHKuO3WTEWroW632Nko4QwnFn8T5
FDTUh9vxee3T24mcXJcb9OtWU9t+2GI7fdsiigVg4dDmc8C2BnsZ7J4zFiXuHqYWrKhCG0ne/AtM
9Dr5+gWarI94tNd++xu4JSQ9ZoXtZybGZXxkM7DKNDAI8IwCyHUT39mbnMyPMN+Hql1ngIKGH1rE
kDql6HLy22NATSZry9ArGJwRWdAtEjKDZK+sbDI+MVO/btSBdDjz630dB49sRYWwsxeuaElasS7q
99XVM9iVUB+e25BpoLK2fUkZYIYS8SdOwwZJoZDgRyzHUE79prYo3sGrs4QFP498PI8JbgR0/Kuh
rWARGdn8VBI4Kq03hJW1glkD/kVAeN3pDpXTqTW62IkbuIeE7io9bFw71OXpsxslZUpbIURssjo6
43qso6DpDUHg8LGLTQeLER2/I7Jh2xGaq7nD3rXM24NNVKj/9iQ6Cv4fiIoGFoo9dQ7O+ohHIfTW
Qyw2BVBQOb2C5r3a14JpXrjjrS1R1KgaiIpQlmwhtuGltx07Zmtbqnj0wl66nKGUxKaxA6SA+GDT
pj0I9IlhCU5w8CQ+c/u4tSiJQZeJdKcfxFJZvird/BxURsR6cpqJ5YjZroIIgb7ePt9Gyj5AdBRN
doj6lvvzHvOJuE89OkCCia5fMKg1zDLfvwCSbD4XClI165nsCk2BMX/4UIrqd/nhV0Nm0jeaJLy0
wc/UqDZDFaeTm+ib480wLhswJEJW8bN8SU0HV7FTxk2RDWc8pnpSNee32V+JHq7J/MjdFnMsN3Ui
P9/JoElskonGfj0nD7mGKac1jxSHIFTYhRuh7todLdJ5oyzKukmw32f7obhZiKENPjIeKRvhVgB3
xlYmqK55TpsjOmMKt/8Nv5Cn6JxNilBRs0rRwPCctc7NW8xym92aUIqP0AbBmbyapP08kIXWxDgV
31yFac0DIqj64nsLQXiLjnOUF4z3k3rUGXGtYqXxR06rpWkOOK1zU7zFucnPnQUMeahd4vbV70jg
+tJMefX2V9m3F2YQ4pxX+eMziKz3oP1SJ8YbVhvM4UokLaV5dUjUJ3q1b36mQ8Hs+11cPiO1xbow
odXNgOFCKfjJVodLSmBSvQsxShz4i6iPIj2I3CTcqVinCj8y10JDEpT5OlRd91gYj/iNxjoP/eJZ
DM0xHNQY8C3Q6n74+Fwl7zx9ZeMMy5kpued0PXeuLP7KgELU4Y+AyRF37BRwLHaFmx+ic0oHJSPz
tvQyXNVwL3f5wMkKeStSh4autF3+YIquHN4pn7Qecz8Qmo2rHR+ADUaDlaRUay0GGcNGjYTpxdy5
mIiuYMCz8uinyqo9FQRY0ebQRnu7p83AALWcw99oZt47erAlq+pakxSjxlzZXWY0WE8WT6vXTsxg
IUmaLgUfMYk5BA/XEohddW6KZjAl7pJwda+Qpc4quD1JCfXytl9arkqhEwWOt8HGT8IwhB/Wq4yk
cfrpNJX2u7aBhwhfmqTPMVQeQa9xrBzACrODspbUrcW7nxR2owtlCVYlxklALyRLi2WF2d04EbxF
Srp3nLXW4D8ju3hkqrDM3h3uAzX3zarjkkH4uxql7I8bQgpKRtLFYzIqcSLC0EuqhMrFibakqgIX
jLJOPPEUS1+hBsF/7hHCFdd5j4mkHwU4OPWMyTK09ksv0qEz/kMIldHWTNHnN96BI2w71WwvTaeK
OI88qgmSedkv+bj0j1l9RR4J2q0Nlpuk3A1u3TEP1aPQDh4qc4jrBE1ZY1Wp4ELnsF2yDsWfBXR/
anHo6jUJ1Yg9trAKcGGdBYe5JgsXWcd5kvlyV6J4prXTbmiayqib7CoVFpPrf+3MxVrxztdsyj3F
zMDNw40ybIMGOJQuIuvmloZq4SJc/M2fk3v6TBMla0ukc7yzXIc54RvP3TEOn5+XujR7KzZlsiBK
3v62NgTzZV3OcOh4zDF3HqHLjrrhCS4ng6iK+pDXPY3IZWGspAeRMPbAW3UA4Ytp4zebObPmUBGE
wIR+mBvYd7F2LQXawNAkoXxGYWpTzgJSsZmf+pgRC7x5HSSP7CzWFf8JEGQRZ+qP/sb25BV+hdUs
aSMml2D2QxJlQSamqFPlepsZi2hMzJXTr51Weabq/PT4rcLHVwE0b/+oGh+jBZkSSQYaB0TZqu8T
MN01Pv84vi6AD/qp4EhcZtl5g+OmnjOZvUcG2GdKp/M1miTvhjjsWQLFkUMRnbSTvnd9nvAzMwE/
YyEVCSMq1nblMLRfCn43d0cU3+ampAzp5zN6m8exKYdpP4lyMCz9r10ruBqmhBgqBzt+kUnZtfI2
mKwGOoFsf4kSkuPLzajUDR/Ub7M2uHJpGgWuARiR0ptCsppVwPlwqzxrxbyROjNgSobxSGekd09E
y6CXcy+xDzZ3vxkGta76fCNt6IWSgxFbkkks88COVjUdR6sRy7Y0MeUtFuJ2csCAti/ZpPoFfa1D
N8Kufeg2xUI7D416iOGCjM+HpcTrLLex1jEjwebdSAqNjXFs/U8jmeqVP2+22Vl8JZVTzffBMrBU
KwliVTQoaLZXdItgn0UXcaL2PMB8fan6UIHo+uknusl7WYB2htQTuy+xC5dRQJf5MjD2uQ2FC/dx
hp1OEvS6QoOLadzp/a1bSraoD6qF5CYBksYHmdukHmUQqCh8Rxnl9p+xqe1vYMMOEIEBJhjFnQpu
LpfBaqGd53c4wxqv7TQOkp995f/+cEK9Xvn8SPcglePMXSH3Xs8OEq8TAEzg3FkBHcrFxQ+TsZxz
QjceMiqzgKhKU4J5Eirckf4fVRr3M38oG7BXM8wAmejjVuzsFOBs1bIePkx8N2CyqJHTvUqOWQQx
2VIr93h7kcLo0Rkw3+erCULI6Y88D7GHEgf1hGZpivdIoq8K5kU3pJRbziSRSRucwcxZzPIp7Qme
p3IcRfQz5TyGMposnr/xdhpLP2XbLl7Zsmo9C+FqvahrHW6M8ytNwBS/WhR09SgEJRmbRImg4q2A
sT5Guen8hyzMr+i1q08+cywr9gz+a8Y4ftq8GdwFkm9BTayENcxz7pdB174FSb8VJ86JJT3XdkI+
fhapoUr3SCNxmmYJrv4bP34znKAe+lDDaIfPW6Hz6eRLT5T/UvF7bcK6B6zA8f+NzWSnpzQ3gwJC
TlnK3griSkEANE0EXMN35aj+AXJ2oUzT5uXEvXPUfWl738LhxMOOz6YC96XaVDI2ZpwGXN1vNCPu
wyj25Spumt/OrRWxkMCxUbNdRKjQ99aIc+3UXwK/oXzO7r0nsZqMUuvfQGvJlLNqLRjeMswaORjk
ogD+HPRpEJ3zQpbrr1icU0a1A3TpKoE8QcoMjiq/kyTU7TJEo4ADqTgXhSDawH4PUJhP9cUk62g1
ch9WyaAptFz5p0+JKogzzj/9xFWF0Vm+rIcqR1m4CXAlnR7MInIXpGm2Xc5IGreMKuiSpRm7I6io
LqI57Da2G8t68MdpIvHD2qCe8ZMykRBba77MCNn8SL6heoDCoCr/WcfL62taDoN7xhqniIFe/jKJ
hw1mrRzvQwUONGFK1sTDcWdlDACftcExguQLTnwpC6s2ONThH1mvwOe2kcTch0I0DG6tgTwfxM78
m13dvzpKQ9CWEsA2ya8xK+8p+6IfzVjpWVN8svA0JW1kI6QvUd0/Pw3lYiZgmf4mycaFhLAs/k82
i2eK5vu6dH8IAajIuzv6xEx0cBLxlalQpPJYky0Cw5us70y8R33oAu1qMbQMYRNsQop/MAekVcIN
kfN/NZXEbzZfo+Pk6hwfLG+Go0+7/FbiXxOi8OKcxYSnEDFZyb7bOZoj0NPmXudqrCzXK5WPRwqp
ngxoBE8IoiKE86VZk/oulWzszEDRtxMSh5+h7UJ3bwU1/NGaIgafeOYkzj/E0gH6b2I90LlB38ml
GFJGkPSSP5NoimWqi7FUzdflebacdz3dbrZApk9z+8gh6NugNRoZkaLDcvnBVMB+T8wjKHkt0hHQ
OZunuONl2PPEe1NOURnnUyitL9SLN1xfTW/VGL+oegbKTf0kSly0ETNrxjDsiq++5mHtJxMx0poD
owL6UNi90X2r7++udotIGswzPkp1eqouR6eIOAyA1l71qbBLyVALB0KD/FH7QxU39sO11iTtxkss
IFJI4SDVhL6hCwoQx0sbWolXoBwBzGl4rUzu2FufMhc2SsE4Bve1B1AnZtCTCDMFGgGo3TuqqGA6
vhhNKSX2IjaWDmqmRPefw/sg3+hBvEu1AOd2182A+6IfgiZ72oPiU0Tvox/5txVkkKa8OoOwwmWv
45zO/T8NkqVUDa+Ilfh/RzzDqT9f/Ybb4Px6oeVCEVGnXWPXCTItMzrle+zmCcaQxlVIKvHzZHfd
NJrc+8174kyoN9ZaH0mBrZsN9Ch89DpWMluk1CitcYjxOiFuY/8LHeege63tA9Kt/sKAV//V9GQI
7e1uLtC/ytn10VyQ3zh+tIXgNO0GZrLMYa30ExpxA2wk3JuhhFfD+2XdoQ05DkWcSTJ8t75ygylr
PENjz0mnO5wb1EK79BEoAmErkGvdvVd9Id3fnUjbObnq4bZSmaBeLdUH65MWBuwYWxnI2PbqNDh/
0Ge+x48fgiSJb+lOXi/Bu8kzhDYZKzW1tsPKnkIWUn8+udHRbdHeqszrken3BSwS8RrczJOfreVH
l4JCI7udPEMC5nrwjmFmvnDUEjJl7q5gNL1c4vRx8OOPMdZw70AS66Bx6ZUZko2GHAbEjrnuzzYz
PEo4sinMokcMXvGFK/MQyeILGfXWikx3J8C9oedzq5rIS1Q+FJIRo+t7oRCS6SmDTFl+wOsf9s9Q
eOdPKr3yGGur7D42wl1kvRgCVL6KhTqScJOHQnij4+eHnqLNVGDquhlqCmYtYV4lffQcos1VlIC6
LD1aliab4PeUyZKnS+yct+gKWT/p1Twgiz7CgvyjFHkCToZ3KOBDUI8rAQTqvKIf6cUOVezk4HuN
HeUoh73HCp6SKxZq1oDfuttB5S3WdE7W7Fm3V/z4eg1VFzjTDpQCEtE1wUoaejopcRVGw66Skufx
OETxF8uk0c6tGrmIyTayuGTfF2LxBc+Hh8zsMOu72dVHszGu5naEBxoWk84AWuaZvp+uMyUkVcJH
eqJVeGl3QSWLyctpUmDkFGgQuzvTpcoRe+QDQz9Er5IA4OSbY8iU0zS4R8uc1rKMR9qOB+6rvqeV
cwfj2UqeBAE2Pdr9WzKfVVFf6wOtBP9EVBEHL+kTMWcJbjFcHB+tw0kdLZuUFG2JwBmy9qyn770o
+72EJblJqGxujaq7L8uSnyCMbO4O3wX8w5hAoTR+rWNdL6MktUNX6sBoqwadqldvHYfcGCR+JDPg
wHt9zPMbEgWdyWmAx4IE7IyGyxogbthMUSA5zklrOQEVZasdtgNAMjQxKKE7HSBdlGaN3P1fKcAg
aS6V/waj55LomWRxgSp1GtW+NejWgEm7ql932HHC85kK5+8ia2Sl/r5tktqE2IB6gSNDNcN4CCjb
12iHC1QF0d0L8Zgd0mPlsLqMCTr39P/lYQYjjgrbCuLICfkGl+4S/BpSWC7ztdQvyPkZ4ez/lysL
dy+ciEpuusN1hZBsisKbdboVdNMBz943u1JvbkZLZ+rsadVrrPYD4bos+N/Vuvlw2vqDiNyU9MEL
3H4D1psJWrh3mewxlZ7E/ChUC0yLTIVYUImtIuqMAi9mjfMdWbWJiAdRrwwM34hj6dmqlth+yiOL
99r/qia5IDpJ/upNTZ3J+/77mfas8VA6AnBvMFcF4CNRpZ6MjTZWJI1z6UWNrX4ac3mxFvbT3fsx
d3uu1azslUOVTlDVclG0wNbPIH6vW9NJtGd/TQlwz4noKXTM6mfYcKJlRKnznEcNDgba1nRcxPHI
9A4nzMGnNJ7vqZZywEITykTMWWAO6drj44FmrHf4vXL8rBbtJWlEV+EAVqhSrxdajX7rimoEE4Lu
/InkVHk+EC359PihVUNb3U8h+9yEBuw3lLPO2oaNmp+gOJQQhxTBXojAuKsoAuwP3Z8yvIrZjGaQ
Zf4Tr8bbrHzoUfCxcUiwC7EVy/6EdB7YcmdCTITi2xiyHa9V4mlO+OzoXnc0Bj7Qh6dXKPG137Ux
yT3Kvy0CmPG9PZwkxxSQx8q6lwQu0QK3TtBarTQYLgwSfLx8i0QDP8xJ8xIVUbWB/m/RbqQTlCcG
dlM3t0HNW0xC5+3IsPrjL9U21mbshm+BgfUNpx1ij4SB2eUp0Mfobrh/N2jyUh4fMSc9/wA+hh+I
ryBi0KsDJENxd25VhkIV+77MzzacSug6/Ti8e5VQNtyd7Y+pNGMU0PdaeZBiye07QSE4tRxk44qy
dfvLS6uMoX+VC+r4iRoi2yTJdnnmSEDj28ERXB3MyfMQ7zaGU7vdVafCJD2z3p8XTno4Ff+u5Bkk
HQtYsFjyDftmpJCLu0WBsDBhy0fOu4cYD0WgUkX96834T8dgdQ6RskddN/NzsqCInU3lOpZvb231
n2pIc1zNINcayRDpHLDHTA0XVR7LM2nTgpd3NRoDnL+eG2hrYGOf0JkX1cKOEowusjVNoFVhD6M9
kx9g6xkD4rDlpAhWU1x2t0o/KFYRo2cTcGkvlKvRRXgPh7YgsDZmqJDEw+Ujfo4v0VX9UwYD2aS7
ueD2JJvVpdEumv4SUedVHcP/X77440dsJvIWjN5uK1ziqmAql0XB8qs5EzNdPn6fb+ZYFVAuqUeo
OQN+i1Gds6+Ng3PzNGUDJsoMYnuSxnONwdG7xy9t4zNXV/O7QasA5r6gMPybVoXZbJxA9ib85z3J
jA5rX34r2mZ581lVhQ1hDCY8Pna/gyhMBrUBqW8H65TTaEzxwxaCYrOYl7a0UJsnAA/oOFGDkMST
L6ei7b3rItV+b0jO4Ai702OsK8o1OEgT4X6xWKGEPF73iFmeGguV9SRnJANSYb30x43uUoY2KYi7
UktpdRUd5lOzhUjorVD25vCXHWA7lYiUGS1ZXhI5C63Z6/J4zbsypcXsH03bBEHt08vf4tCmuxzY
2MQS+vtbM6MC9edv8vlW9g8XfRzK31qLxAs8qbd2pLEP2oI3x+qDXrGdvVoHd5C4ClTKU04jzb5N
+Pb2GndU6JtotuoMV1ZFctNp4LCXMDlwFXXM35zIOBq318t9FMdMVwIG/Sx/gxUHo79C//Mt7dev
/oAgkNiYarKY+yNV7bYFUgG/v50h3TsefOsjMebZtglhJDjxlYyeNJUJ+qyTUCjHrVmVtXt7jwJe
DCTkJhTkvxjIKYcH+jCFytz7YJzP+5W2UGu3HsE7esmtvLHR3LBm6rX49+lYRQ2+IE2q1Rx0rvxJ
jy1+5SkEBZjoQcxVpwLkdgfBL22jGiFmZxp5ZEW0NdMoTBIq5Z8rz7MEAuCwiXVTwMbDt0KbDp+g
T4XSCKkKlB/LZKL3KDYWGQZzvrjOd4SHL42ibhgj10NwybdU9yxXsGAmoT7MpP5ljnBS3+T3ncSG
h9IkTDYxP2H42/tj5O/G0UMgS58uLEhCZJb3X8xOMks1Gr5hv1mVgtEYcVd2e7LBbZz0cf8sqN3C
C/vcYeIC3Q76UI0hYSNirrXEhhBY/RFckBDaL0BJ1D7wwkU/RzU7qvqFHWAsXeD1Hm/Sj2ajpYoo
Ec8sEwVTzybJdg/AkyyDgjMi0bcG8GUYm9rS91GMxDAy6QHmhgWngsxWKrAog1Ije5g5hbVQy+uf
gqZLsxtdTZbIpCTzohKobJGNPRN00aU8R/nZqaPXaJgtSfLTBFBVZyqJdE5/2JofD63IQj0n5i+/
jravl4X47AXgEILEYdU0Z8yOXhRMXWTRfzCV+lJAp7n7pHDUGshWA2atf8agzTCy6vZubXkLauTb
hPh/pKjsVN7ww7Ax4nsaFpEFc+lpOIeDz8mTrVxvJ8NqR6wo2siIhEGOiZlFQcfgrQO6Ka9wD9A2
GwUGqWgoUZqi3JwfHWjOyZyiPICo8y1/kZNsKGWXEQdPmKgi8lnTFvp6CyW0/FgwUudCB9GVmLKK
jrGKiEnLs7h+6bQpey/gAbaltBXgy8ZcylkVVEgtNz3wB/w4PNrjAltU1ONXpE2+n/nBAlO1wR9B
hIKQ7FkDp+oUy2P31YpUX4UFvDXBIjlocTYpBbZ1ibAXPykzWJTuWf3ivh7fOfw/SjeAjVqmBIZh
QLkB3+/nNUNem8RTren2eMTeiGr4xsVZIC2kklX+sFbKlhoS9hxFIbHHsTJ9EvCZclg8wSxNxqWd
Z4bnwZK+qL7QQs0S3yZFHj5NLRRsq9nnGxcVDIqQUNAqSZ69Sp27GdPQ2af1gSGlzaZtpastc8Lh
GUlodlge3v8Kj7WHnpFwCUBgMXAnQV14VvNOfMMSlpkDUWMr/7vRQXrC8JjqROx0Ja797LpS+ctF
tPrJVKDfnbguN2d6BfSsw16QqorYcbe4+FZINFI77q76fmfrCHCDem0AtED6hPLzbECnFNCvsJSx
lzEEmfudrXn/bMbZIJZXz+iEECYS3TEsX6CyXrKcs+3KtzBIQ//vqferpACn6q++v7UB9j/eFWTN
Q/jio8UgCpBgqmcIspL8Z6o9X0t6ww6P8fNKdLLyXvhy3/vIrUcIEXG9DJpiNwkyElHp1gkxSYVr
xPuiQCHXm9Zhwcxafbk3fyeCCv8h62WaUhQoxMEUf6x8UFZgHvYJMbZr+usflfoaMpXW5nHFF9MA
m/vnZsg4ALpvbDev27df3RNdM5szPqojEwQg3iMUsrWKONyRt4wyoOS62Q1g8YcO5MbMAINuP1z1
hNf6rwEWftnbQJW61WJaZPH2t7i5qQ9ZOfNcByztj6yJY+IG8y7IF56HOeXPEkRQcHWHmu+rb9Uc
JGOfEXoSgbE2vdQqy4MBT5XycH6tt6tiZ4d4Dk2C8SWcpLSYLW08k1BwxKYd3OP0vwkYWog5l++F
/Y6Gi6MFbi5vGvhLm0ImSbbfUH0AeKKoB6nNKT4e8obvl1EKXLkgr5Wgi/Kobfd8n+Sa039LN8yr
AFuq/EjgwKEUv8MyNm1mY3rLU9A9snIrGncfIpa62DrOOkhL3I5kU5lt7/R+WrQTzEoYiMUPqxe6
uyA2IMkXTZPOorTZ1WiGp1UekCSYXMogD6FZmlH3vbe57YVwUG25VAIeLVwQ4Dt9N4AMsfyuLlP7
IZP0O9JhpYj7KfMtsTjHv5d7IfA04dRVYhX+z6bDfrFPPjPl1AChpS+ihCeAXtCPFtGq87CQaAZ7
ajKRv7cIYoHRNMpddA1JToF2LONvs5A/wyAeVMafXXoBQPa2FbDFCuekcAfkPgKefsDm5We8W8ID
UwMOQBgXweB26vrnUYBTcodKYHVTAyApukSuzGNs6LMBmwIrcRBM/LCsYHJvjptPJh9hgAP0wqrv
eehqZ5xzimAgtM2e3fFQXPKbxMYG96tiGvrP8ATi61VSEn1nsx4wmX4QEhugW4ZttmXCo6e9g8NA
2x5QcVH2lJTHentZpJL62AiSnmflTJtCGcd8bCEsQKDqZaOXeE7xqYg1hvZP+CVv7wvDXLszjbuU
gMcAW6MU5yXXhF4bKhQzOaJmVMKzXXtOSD4KR1DypaGkL5nM1QDZdvv0fc1hDrwM+4eZbvfQJxEN
2KXpQ9vn4L3rgl6kvj5OINrXmfGhwEaocjLPknVItIKX/MfXlx6IXBHorMZLD2s0kIj79c0vRTAt
sR4yW7KZhuhvZkDIOuBsW0AYMjiVgSpyhE13Jy2dGU/9CZ/4RTxKlyBmOFEfEIXSsGF8xJezcSjF
cRySGssjFLY4d8rP9EnBd6ZUTXwZe68GKXYUpTuy5rdFyYRbexS0xvNF7JM/ZqIwvvq76zfUVaHg
ybcdMvU4HFYPkNQ38N9wlGcjN5km/nbRUxSltsA+2pyOEdaHE4ax07ADbqy+NYX6BaVRnOrbFHCx
q5+5RQzmbeCmhR6r1TDF91dyCJP2FvAjciP0KhUysYUQiUBOPvd95k8xATFj9IjHuRIe2gdkh3lG
7dApSjGmP5Ix4MyYUncIxUysvjaAhOOFdSnEBp0sIUiv5KRT1Wjr7qwJWj7n8NrD1wgndIKGpgLt
4JSbSOFGiqdpAXa3REcoSjflCwRQdA0/SMS8lkGeVC1a5TsgPeOHWvobvvgFAnt3Z55S6m3sdgbU
CA7DQzk0NMlNKgNLwnCN92tRbny/gaIYGsHIpC58NG/EF5dNwv5cjv9wdMRxmp7DrGI30hZXwCUf
mPioopVTqBvqXM2w6mfJobhbQm7oD/LMWmIoSAZgEufQU38bwPCcI37yYqVJAHR2MZqtoyU5PjWR
kA1XB+yM8reRQorJw2Fyceqi2XPPyJipjZK+376M3j8sZQzd0OklhkhlPezDmUgl8emruR9Pt6GF
5ImXkeZEifwMphz6HHAtD0rhmMzcCcJEprkTEZYXLRU+s/2tSYnPmo43DJgC4samtJzSCfZeD8X2
3AdUmUzG/z8kp+YVFlOn6ZEOWdsCIntPhTvYAu/EY3G1EkCIVlBz0o3ZTAPS7Ak0BZYaXelSe9fk
ySFEH2auR6QgwTPBbeIeRbwu9JdiKgbSD76xLzD3yJifScMa1wChrwS1uHawtx5qkS+B76Y5MuV5
sLOaXeQjWskhy2Y/l2d0L+znbLOVNSR3vnMi7y7OXJy1Q1WeHktwn+oA7R+0DQEc81eGtUjiHRLX
klzbix3JC6i0b/Mp/mdTtIQaP9G1AIAVvTVFqbzdGRX4NZxXwPyCTPj6N+J3Nxigxqf9oB68s/TP
jwiFhTCxMMpo2gJVtYQcaNlQtaajI8aRs5060Nx5jb52wk+9ZJOsZWr4mEL+7fpRf8YFseyTEwFT
zicseO4OXLdilPqs7mcba2QHRVz1w4XCwhGGsdQZFFucGIYOohWuVlSlJ/+UF5YDEc5uw7e04Ndl
UEr7NM6vrvP3lwq6AjzvwSdMKnlwUjjx71vXXXDdxEPLJ21jPkouv9cROcOvQ+5qWbnqQxcUy385
E8+WEA9aZCjxAWy81GGldsEAjqelAvQsfib1FY0GtVobjz5D6iHSU84vYCqURJqwZ6YPXrN3XEV/
RkvOL4fvVPvdDzCJHfeZh62uvjgvvcJhQ+8EFtA2Y5x7JXGqBSxM+rJbaX3OLDCH3S8PA6vLLj0+
+jHZ5f6Fez7cW9N7xwHKmaA7UIis5OO7iQXXfDtzUhquphluf0yhPdyIDrDw8SbSULvKjx0YHDh0
wUQTqhdSEYkWf/iTAP3QtuqiIYre+wAgrjYUXcKmeUl+4F17hOuru1+frkDd3mUtUXg3kh12FS8m
EcmeQUVPvke1v4xOp3IuHXb7lz8jmI6aA54ArAFv7/IMjYVkcHjRj/rAovpIAb3xNLRtd/6dYCW9
l4brR+RCcm7dSAkqL5GaJslwAxtdDewSlUN++fLV82IskKyDTkSN2kLbshmw8wGx3ohfvpTCi4JV
jU2at+wbTZ7m/w01MSOjANQyWTJTYRlSryaj3w2m85RWKpAW+/XmNy7KeKuRx6rD9jUNGgRTiX8i
Suln/4wvngSJSRfBanDtPPpAgg9lOCWeicARBfc01eagW57fzFc219ApXc8qqIcRyzqJiZsCe8NK
nwkkCjUQcV985a5iT1Eh/KJFQQZWqtMPNYGNpgmWqx0S43YRLQBitoHDWEtSOZAYqD5saaDix1OL
peYed587c2wc8cdkc0UmrKL7Z0IqCpYixVqm5YXz7aFkfML+SQmq+9sLHgpoBDKYADp5F/fN1bdA
/yayrdQ0HuGum2dYcw02BkVE/LeVOCFdDST07ppCdU1hJpm/y6QjR0tX5LKInOCc2Lsr4nZbsvRH
MQ8MixJUK5xmGeWYMJPNC01y0CYQwKhTHzDxHpYgwlMQEJoBDVY7SrAqwalzzZTKZ3VaAT92rjMC
lIM62/dQHztdqyxJXNEgqWH19DHYUcR/xTzVU9ZVYeGlKHpZ+JIKVo77g1NVyWBfaJY98Koime1Y
Lzj08UJYX5q4ngLRdOmiHsvufElnNQ1iaVZ0ezeGUKY3GxEOjQt7CclCfKnqZp6ayzQMZBnjQdR1
Yftinvuo1geX3heJF1h1oCfgSQ10qHBHFMa0Se8jNUBPY/p5FV/xbS/f0mDe+KMFVozwi1LTGOTY
ukFx3z2CNO6q1SAgMSYJwLDXmGlEM/GVj8/FyzobxRnJBrjwB65lSXrYlhYsYgt+keaR1cUjnZ4O
tmUT6eGqvFvoStvEDL6oD00f07j/cE1uoGxDuOBSOeQxN1ZdNOSRlx37dLEMLngAH9MK21Uh5XLE
fPJwLd+rJgJH6RAEUTDZ44RJ5d56qNEVX8SppzhsQw4gKUX191jNIk0OioBw/IIUv13wikcQereC
GDXPiYpHCK9TquZA+TBHuTlAHiYyGbsU/Th5MlQBfW0+9OG+BDsWtmafyIJRuOjlNoTogTrs2wqL
28n2BdoPDJvZYJZBPTLf3xjRqzPkpFXUFol3pZJLg475dD79rSVB4685uuZSgHR+0UDVouRuXQWn
g8yMOQnElXDGYXwlzuqW9Trd4mF5fCTOWofjMehO3uerSiXqCVOHZnMPaJuXwsPp7QAshwH/hYme
/XTy6f4A/E15isK8mpwQEdr5Z4kD8B39TScXJn7oUh0ZMGsZkk7BN3d4gr2qSxLolhRwrIJOpina
PyzxAlYIedbeTpZln/FKw2p7O/TzqnqcUZYAOkzaNZYHSkOwL1Lcz4fkhaqr+50Ir/NEn5kYXZTM
I5CW9ujad3bWjYhSp1xzV21fqWyHoi8uEHKdlska5+Kr6XkVlLIyqWqX/P7Gqzy6c6PKgH0D7uJY
WxTih8QALyFY3bkYfoLC4X0pnAEn+3t9xu2NRUO/1vgSojTRweyw3r+4UwwCgmbEG14izgt6uSXp
ekkLtYSTq5LoxPIo16jby10zYq4/pIPDRs4r4zsUNiPf+Ax+v/m9XB0dF1zL/RZ4BDYfsaGdNtwJ
GVBFeFlZku3lHy6P08eZJjw51DsTRpV6ToXFi2tBPeD9Bn3HAeFZAaxqWRVRUZEH5ERT8C6R7lG7
rMZeYIs+NpOVGAg3acxI0bHB7Qu8eGi1oCDXwdsPjViY5ChcshXBTsUuX6svw1byXI9WPa69xl0/
RSeZFZxK0gKrD4usZft5SRy/+0zPK5oiTs26WIN4lpe28rGHVkgniZHzpMoKFqY1zWHIWhqxbmGX
tPVOtSFVmKY+6hMZ8IKak1Ltp2N6xOF7ohsItQKMZUw3iM/x170Nrg/+dIS3sj6/ADVQEuEX9FK7
smowpzNzW2s+T4WeSRlbgFLKdh83GvjGEWuAu8WH9Nk2gzBnr86pR+C4HxsYY5I+QYr+9zOWX1T3
ln67Z8EWUTjlzMMDKL5bvhBrKcGSmQLGMR9QSwqAUrADBclWd1VD8QHI9zsIbpw7Ax/NremZEgzL
IUb4t3k6Bi/wO16wCBXGqHLFealf4X6XHx90bzKSrLynvmDL5hJj8wXcgltPrfEVER9OO5LKd1ad
h7IpiCD4Alv9XHlAp5C+n8gwPqL8w3hj4vBOdXa1rVuLhcJjXKMzllIIP+NG08mvx8StfNMGNySy
w/3JC+hwPPA5xlcBE3EzDQsGNJiNK3NP6sG/DQmrpV0bx8dIJegGwjnsQ0ywWW6AIyu3+cDI9VLg
Pskl4NTW40sJZza7pHLoCktXEJeGAMPd23iG/AgtHxdwnISn1j0SSNYl+ER1WgVFIMY1nwfFPsFM
flIiHAjjHXU3wX64JHO+mFc2JEdZb8Oo/QnRgG9fgY8tbPxU2LyZJZ2w6Qtt2/WZTzL/OWjkVqYV
BaWKRMWB2YzluwwXDgXnqTO28T0o31CCk4CKEkD+WfQ18UdVRExBalxaGwdWYxXeXPoJgEhtGtoA
rp1m0baJDY3MTQfu7hYHYBzfFWLYd/WMbT7V0sOan4kYXxMKCpXNdVsavN1Rfeoekym/xAu3/Za5
WqYuZ0WWEIKD3Dyg6+UG97OudlqVSa2e5wxeFe/WmbW9D6nfkZKa/dEviqjziEyGtmASYq1ydsVb
lkawLe3lExVoP8wEIRabgDnCZgFcu03gXDeJkWY6nGawWLHvlt8LcLtfydD9idWjD92hfHgx6BHQ
JLYdgjTnEs3/oD6C4eyFX24z3Ty6/CfGi1jPrh7xz5cUkxE3WU8ZLqL48bFBSMxKagXzIE2xon/z
EwcjmlE3QaQpZEACikwUUPj6WbU6qvANT3ZaSIf5vj3PjxCdNWwaVMkXrtrQnVtg5/GnEEwgywWQ
4p9zMAxzVmz9x3Am97Q1Tmszu877qwtBHApNAPzcpNivwux4f9xweAJOvRREMZ7K6/W2nLzMDg0U
nBH/nqs9pr08Ctp/E3Wuuf00YoN3pXjlpNTisOvZesu1cRtfo4PzhzigXaETghNJR/oJKftS0Cn+
DXMf1IKbKNmp+bUslgzqpZFLLN3XB+zJSKuQIdwA7Qp9+ZMwWCSLBR5l8nNDa8vbI8v0D8mnmzKD
b4P1qilloYQE40kUABgPRpDK4z1KQEkXQFSrg0YfIDxFEZbQYOIH2Lvm+hWByuCkg1hV4nT5unGF
dB2zi+yprKoFQXEXETSKOddkx4qGQj9w0lOx29Tm9FqAwVhGW8JWjK3oQvnJE07AozySN4VRkCil
ZRTk/9thVsMY+7Yx3cD9RmFMCv0tFUao5r9TQkKu8YeA2j6iZGQfSGqi+Gf+CIFM7k1y0Ytei9+T
ZHL6RZCiE6vNzMP8qhFS6sd8+2GoAV3tDQISAoulzmQQR//7zZe3YaI6W8okNB5u065wRJdYSD19
YOIKWymH/dNThOLdfVeTtnFXN8VCLgm4sP8EnD/xVR9Mn914yRXafYQR3QtXPnjB8Qwlx2FVn0Ac
e9v3SXfOuQoIMvT0KBxeRv8GHcpsCwvDui3qq7TL3OrLg0S3S1fg247GFX6XSgVDfmb1RI7XiUSh
rOzcevqXNMJ3pVglfou11z1Ya/QEOKoPmBv2+0ZzQIx6/nrPnM1xcbxeWCNX9BhrFAG8oPTzpg9N
kFsVFw5um0spxksvBLbZNNk4nx+0KPQkyIS+xtE3ANOm78CuUof92YpDQIYV5MghBcr0A28KOisz
NN62kIK+LWplF1040sSRTUkIAfpEb/k6EYZf/0mtPviC08VON6EjNjhzSlCvxezBMhfzkd0fZoqj
kwQZNEXkU4pDIus9yEVdNXPDfS7quvnBUbg9P5CHQNatUmf6AowsuLBOxcU2YmGJecOqLtJlzWOO
K74b5nbHpsxIvb2BMEoHErPFP3Pe5OtBprxA7GCCZpM7ckLlts2uWJ8mihlARKZTMeHXOMdaC76v
gRCqe3moTNmACPLih6cz/BIt4vl9UqjZP4JrslkUmxeP5p0b2JNidzroBrKpZ6RklTySkTLR61gZ
auMS8wKQfIha4MfeSxSkZ7Oe4w5i2+qVFO8HBOiVCO2m+L+xzKd3pghZlX+uFNZ2uMynKFPumiNt
cnutqWuffCZpsjCOOc3V5qkIrxmAsHuoRj/ZIILdYH0Nst98PSKp2XUBJgkHvYnStHeuIHnrCZUF
tnTWs6JbgOWfMJxRRdDu74bPBYssYmaLYqbIfE7DY7WPkl56r5No9Mg4h9FzcEnXlYEb5Cw0ToXt
D5jbmQi+aGQlVTaP3sy/KogWWXJFbPcmjsd6kCDsnAx3ckImC/QozmtFNJuV02U1qoqNNTVihdnL
ktEEMODV74YM1eSlsjE3EUSEp0wsCcfKzQPfUD/LGopHPYHc0rvDdUYJObrmOAd1Xq+gk8E473FU
83QagT7nTA3zwYbhyp7fI3BwelXtAKdryIX9a53Iw5zeMsj8e64VDbYJ5QHROJ5tpwMoEkwTttjV
L/Tx/48J2wcue/q4mAoRLBZCIf/RddG0qSQgii/apYA9bj2vZpT25KhwevupUl4laQQvqnO5leU6
S8akgDGBT7WVUh0SzT+sdTWhz5AwV44tTjCI2Xzbqr4Pc6h6lqPj1HUuPP28FY7qu0LzC3mePkYs
CBYeOKSUsqv0BStd3nAqOc4lNLHCgmXyBQFuj7JHwEqovSUr3FEa0dnk8w7oQQyyWexMwZKhWxZH
KbkqwJiwCoC4uWGkFoGuATOmwoZZ12y/DETJZqGaGOzyNK7NGE5y3KwueSDkyQcDGXawCeudtV10
gtxu9z61+aAydZTNEPLQOz3M2zZ6LWmNr/LAYEs2LHI2y0Ua0NvhuGBAKAfkoxoZq1qeyvt+Omcy
gef8c0yietLmbOXkVveQhjLv7BZoAWmWDbJkrhHND2we5Bt+ho8OKySORWylXCWUJ+vndZzWOed2
JwXgiaCR/zvNbrZ+ZQ9W0MOAwZTSgTnTK1sXxQEfybJqGNPUIRWvCcPYznbNCaxDyB3qbz7KpYqv
ZzFEy6JxGiagtBvxxJRHbEt6UryK0eVfpJhD3JrDnRcgnsMP+fQvx4EhQGw52KxWVcum8CHffhhp
rOqb053SdnH0q8ijSOYFXXBWY5U2j4YBAmhL3p7evKZztS4dnlN8p/J3S71fIy0r9cGgFAgAALr6
2TwdquDbNbknU2xMjwPCscTy8tS7eq2CZ15tQM2f66uJAWOpH4BCw7LolklecRaEAmRHlf7p1MS5
3oJp5P+z2xh3YBwc6kFnpUe5mreVabXsR6bIQq9A0bvxcrG4as3j2pGYZfqBRLr62uO5s19nFTga
ZHnw5swGfz0gLKaB0fMbtgkTG3qVQzXNG7gVywyuh397+nRr2N1X49u/SXvt1SHCZeme5Lr2jZ8K
ttUpqDQjt+pCE5Jlyn+gj4Xr6bh6L/19jGExNuu6iUA9UojcfVUccjDAgsXjV1drQxqlEw/35dYI
UBwJk663iKvRgouG8Fm77AgCrtJuCVCNmLTVi/6Q4jbRqgBR9EbiQbBiCKVhXSaL73dWzvqLG6Nn
qvP/Y9A3GXT49ElJdAKlaxo5QBrJA4I1kyY9/QsUYVx4cjPthhXdpLAmyOsO0DT3mfWCnxSehVPv
hfacdJsXgAYn7wfGvWD3rLq1VCBeDxrQ39TpKJUlY2EltEjpKHuDurxieLLzO3q6fq8c6Y6Vfu6V
3xToshj+gKyDdw/2a3Elb9aIraeIz7dSLn9YV2OOF3yR5UyJbqIn8lkJAjroFyWq9waM4tuNjPnR
l/zrcU7Wm2F640NkeQSDu04jgxmld3MpvEWNooZbxup0pDg2BfFq/pJbVkFSBtIdYCBrWVpyyNbL
1YgxFWYDz/50rgQ2WVNBTdv3fUxVTCifAVynHmgn6LYHbBU6ULzK+Ix+SpPVmo8xtzmFG5fKsgHz
asc6U8GNJ9YCLRqlmc7Vgb7quuewnY8D5zyhHQ23EvGok8gOjpmrAi6/47Wqo+L2+ego9BI7odhk
AWGGa/fxrdNvJilS7O3vXxGvIdOHNXHq81kjfGcqvmeDjQJvvGaiJ4wM5O0la7wR2Ti7tpmmNUup
aHhUV5/0DjJQiUmdPaCJpFkBk8LA4kqZ7dyl1+6nIUGXxQe9/AHOw8CE+naDztHD5dwbUWyJiQi+
ZLVkPanJt3B16HjF8k5UvNgjrAvqBNylrh5JShcjy2Ta6hfUDGjBvPtal/5yGyuP3TaS2hsbsrnJ
jmBgtgpayAKGLSJbSMwFv9O87dOBlr+uqpD4XzjTNJtrN6SEKtkDWdLCu5ZpUEDtPr9A45sh8WjQ
dz25heL4YcoNSGnRoJW+cs00uASqaL5sSqpzls+l1nQl4RtTAOcNtbH4ap28WpnRy4znIJx15V6K
sjbMblVRiNJN179p+Ux3hIxhNPBts0HluI7/LITr/La+JQKPfhZmGHsfkhUrdB2wQDCX/753Kpw3
95d10Nmf0JLmo0r1/37Y+ozO6irnBtwLEfcsRLQsRfu05G40nyQTxobK9QypL9DyrMobCa3BIzWc
X3Ma7Aw39Mwp9pzhNkuWkcG60D4TOaK50nN7wOwKUh0Ehz64YbwXdOyX0P0BLp38J/g+qAw1Kd0y
BlXrEL8q2SgxyLckDSktqrS6ij7Ebo25ce2ZmhbERsTKxH5FhaWbGswZiBRtoyGBLz/Mu0Zjqurb
Xazc0bSmnMYHQxrQMYC8fNz0setiW7/GoTDwdWdn1tp/y87MTBXixfswdcTdgCcuxiWjM+910zbg
9MnJV9U8zAF8Y4EPkuLTPs54zfj463B2c8jKRbl55eN5Of4trrG2ekHy88Bk7C+tIVMlEV8BNGJK
Hh/fCi+Eb43VogrVQChVCtdo7x/p/Gw8r60Qmd83bklr4xCm7X/LD5wChDX/6JqRl68Zfyh+g0B/
SRFe8ZJU+UwEUVuVUXW93Oo9GMSVbp0KEHYBUtdGvjl2Cv/nSTOfT8UCdTJH/eZY25EGtk3Oi2Ev
Oj02qYbfI15W2vD4NhU0vaOn61TvfABlobl5SC8AJS9dIwWWd2qTl37HCUXtxFHJlnhi3l/E/EOv
BXF72wp42to20XQSQX8QAA7z6dKBR146lvF4u4BsXdtCFuhZWkr26iH2EbZopt1XeRFB2iYWkDIS
/xVcmYzeMVnTv83uSUrcgefg8sxjRlMc5dnWEmaZ1SmfMs1gB/0Chf1VOW9ehM4NVT4qKbUHzOme
2MjcsiWGZaa7xQAbvsUZp+Ix7GAy9w5yYy8gsdXhSY4qi0fHC/dAY0DRNCpipfzrURE+q8U551aJ
9aqoFi5EweZOogTapXk42+SH0M/b16ePSTFDK4AqCkalzqQA9903FtgtBgfJg+4SxX8bCNGTVGyl
loEupMB9QR0i7Hr5gysu8wOCbhU2lQGzjVM28tyyJPifwcrmNxh7bc4xTn+3qoGUlueiiUCkh2FV
iFQgYXFtQt8EubOEbt7j4hQ2Q9eEhEWbWgurkVyzDK9Rb1r3wMOIKxapKHiLINETcMt37bIMdseu
DckxMjH0YG05/XKs4cMd2FMWOYP/RIUSwbZoyU6hb/ynq+rW697DKZ7qKy3HT3XtHBFpaHc2HaE4
WhVG3lDQ/oD6w/uJLwrCBrVsQdmiRUKVl/DG5lFNUpBbhIm0LchpHboFalKIvok8RYWquj/T7RAL
deL0uZWWvvQhQ/nkBmhVfhBI9OI/t/+KdMqB7JmDN4DBVp8mGm656Psst5kzm53nNiT7vP62avKC
cQLPcCliYrqG4MStdTaKkSaiFG0mHlr2Jd88tXIP5OsIggf0OeXsl59PVyzdCkJhjiv1IsgSK6Hr
Rq6G64ujSXvlGCYpzuCcGw10CVPtuI5itRJAi+Yigey5ukEbUm21tZBy35GvIDCcV3flkfnZWW9V
XblMTWfT2GMJJB6gtn+XDjgcfEzKBhjat140lH4nCYcIcLKBMQzOzEHyMyVOb8XRmd8TtDfQSRb1
QSOhEsz3w1bYTmII8gArT9rlrkfIf5tTYWdZlhLGbhwnJP6WSyj6zrk0RzvO+jQK2Wf2GDkzvJJ3
iUDFaCsYYyRMwVS9bKgBDHNe1L4cUKMBY9uWh8SpdQ7oXgETOJuUQMFXUn+efr2qy2/17PPTIeeN
ewLDlpRNoLe+vXqPhg0DHsNXKORZxJJ7KlUdGyp+Bj4thLru9LaNO9m1hkFzGbqi6ORNwWRVdioH
vcwc/WSk+puHdkiKAuWKB1iBtWACK+x6o+vk5xavk5L6u7xTqdmKp1DglHojpBp+riowEjomx8lo
uF1Dd4M9oSwvrn5SkOFn8HOqnLDgcf1k9SfDfVhxkbRE0ODkRiT4lxUPssS5Yhi2f9029TlChgzC
WSUeXmKpVu5JoVs8hx0bDU2GojbeUMk/bnIcw0MVayQbwFmLcjTq7MI/NZ1/TzsHXIXOW24tqPzY
9Yu1UuIfQ72I/tFPCN7VxFj80hTgcTJhDUOlFlDvaWPq4pGFxoYNkefljMT6fChGC2XnZZuNFoww
cHDn1O4yGgdm+OldzAfbzAUD2qTuigF0/LOUy/gAayYYBlq/dqWb2jNubobNzueWj7VwaO0ShJ/3
LSRuEjcLrgEnsLAfnZXbG9Q+H014bPXVQwwcA5qZDoddNRxgxjy48pBGpD6bp2DmEZw9XqJDCruk
KtoqINl0MFVGNpoytn4Jn26bQ1cq6MISPGixfQ3yAG+SdHAsPXdct5HiUR64IWyjNFzCoOi86crT
0DB0TR6CinH4Jbj2I/zU6Dt41pCysUHIwU8S3/Rv4mknc6sJCPHYMFS23ZJFWY3dBYcrEfOhmKg8
DKfB2aX+3JqZR8PV/q9a01HQ5gmTBcmMcE7NZeZbKxQ6pdlYEeNwsT+HIftsfHLBL4tnOnE9jE2y
slOV+czqexmWzmQGyacb9nkVsfBczcXXmJiDG9AAN4RGIkpWnPrq6wDU+XmbJkgLfVn68t/B1Jfj
NesDPD8h08CxXU2paHCx2Gn3pqIWId/UFUc09usRuiVkgWLPp8verSVF57HNHzhc8SkzhGw8X97d
+k6L2s8ejqlfHNT6KtF4oEyPDlwW70mzq5cTfVbn1y4U0UYYDVOIiSlqflZZMvXtlhBPZkdSsomn
T66gP6sAsIFsdU8LCYv0sQC0FDm+ZliBHs9m3HQ3wYtRYPQ9s2XmklxTDQu6R61GiN+PtlQt1h0P
8NyPAyo5qu0xXFvoOmkhJtAUJHmejbGEy1kUYHi9jdsEBCpAelf6QP+Lva21mBtAZ1NYJ5XEXoJX
BqaI+j6oPuIspPVrAUS7az15bDFko7vOYE6zAChFkrXw++DkOFowoLpOtY7n/uvCMeysVsRQWtBe
gpNf97YGFA4HfYbrNGOoI5bf/KOQ6QcRI0EKYf4SKaZ85fVwgxP8VKDoXvMqKwPbQVFtjasulmdO
f/bl7d/xgvT2CcHEEMJfJ/IY1rq8ydbYLbQK0JhorrmbIhS0v6/4g3K6JE8fHvRvs+cYOoX7cyAO
/gsb5sbUKj78l1LYkZdn6MAspkKOZSqGUFqsp9Dud2wqRoVRN6lIWXJCCYuJSUGGuq9TQLhVchkP
OOjM4bKfVDyBBejLECCaV7evezvz47rq6bFGkXwCgbx4Wf4KOCbENywOuf9Jn0fGUuGTnQ/JWJFv
ToKlhv7vNPUeR/72+aqlboU/WyP40Ze0AQ1Xwg0kYLDmCBM2wf1c1ZM1tqVNNdKry6+WDa+EztqC
v/JEkCLeBCGLRP1NB8MMvG/V+3nmd3i2bP5W4MBuYgWUZS7vMTA3pDB6HxdjnJJruB1q/8p38zMV
MpoBFMWMVTDRmtsDKrZ7FUeEtdTnAQWV3XTHmxAhsFOX1BbAuyxi6axHSQCDPFfZqqhcAyS53IXN
yVRWU8oVhESLYH4zgvm1cxOPKST/a5SL7FZbUF0b1NZ1mnIiDhjeS3dYkqCxBDA21SYiUtelX6rQ
SDIb5FgrBnxVCcufox0ygpkGulzS53rKmPMQ4isuNKjqhWhWdpF4q0hnXLB1u/vpkblaW0058vPN
DDCm1yQWKglmHcEN1xvrGHHdpyOc/R1uUCO0AHMC8lHw72aLh+p1cV0QC99nUG5bPdfj5vLwQika
RATHCaMzT5kMSBU4nSp5tC3eOoR/YNrH7oe7I86zbDUTj3abRhGhqSdwI2p3zCBjs6K9hBE0CPml
UF5yOxG5tfyMtiMaD0CViP8u/w2kMQ8PV8Fpw0QARBq8KKw7oZX9ytSMrcOcYNpE3UerMuF2jYFT
u6IQov8OZWEKBD4S/HtzpQuHxBXaP8CqREs88kRt3L9XbWSk66n8GW8BtAhp8lOa618W7ElGw6kD
QAXs1Xe+tk3+d0mywyu2vGPmoUZc28eU23tCGZEOfCFUyb2qhVpH4Vzd6pqk2cCYTIKvo3rSu+kd
GaByq7xSYobG9t671Hp76Mw1tgD/Q9F4pSDMAVXoWJZw7UPwsGQI2t+yzfmJxOXKCiBFoFCBAMMM
zkrLwiKxz471aOH0bC65IEaQ7NOEEC3YHaVJsED4jKKTwPX0jvR+z8YKjneaY6EfL93wY34zFdUF
x4gwr2059kqxr4KI0tgSzhrrtfDfLY9BUy+OIXXa3NnthZhR6a3lMxjMvP3QylbbH7mZG5hGD9Fl
AR1msdkTH6FyEUyn+6+c0BHb/vy0nzAiOiF7hT6RonvF1bWxq2KJEiikxWjJ0THemBdtrEoGXw3I
pVscDK82IhYHBMS5Te9eJIKpFSir5Z/lYd4VPKfpQw40+A308Lc2ylOl5qIn1qjtdmUU2cYqO+nx
zrtgP1MsxjgU78G9F2KuiPukvsc1hGLj+8hR9UOXtcXDNozudAO7YXe8TYHnHVc8afeGngC4HAop
NaCMPSWMbu1bzvGA6MevrH3KXOzXmuAbgXDgiD8pJhPifpgCqUU2GGkVvEy9kBtDuObiHq5oXrFy
UJJw22kMrTysiYDesoHn+Ds4iiRqvM4NGj10fZGP/o80ptOoVLizEKpGHT+RzL8sgawA9MyjTP1+
VP+Wz8yT7yQMEtOUnAGLgpqfK/1kQSKI8fS/EMO181UKqxkmlNol2MP86NtIQbVY6rYLpbTkWhoA
36QtcFmdxmsBpAT3ildzkbur6SZp3Hys+Plyw+kz3Q3Ffiprhui9icbgGyBj6dx8S6pPlg14M3y+
dlV7+5EiPGQfNw0BRGa4zR4lgBYX3lIsPMRyK36Unmiijo6DZd7aJweIDJugvHroybxS3N4iXEu2
OAJI5z8l3odUWjGE9/zSp/AyurDwcTsSgYP6i82rMfrt48a4B8ODaFeGTaCUKeEoU7tjPGPHAmtl
OCtiPHKKqinFFoVOScKsVa1KJytsyKtdgcezR2R2gUUviZL5a7USDtVVKfVrhN0HTtdxLitBxU5E
XoCnZsJGn1+/JdTHlVNta4NVvTKdHHd/jKH2EjkbsX081TjzUZK8hK0Nvl8dNViFwOY52aGVhWr6
91xfslgeKed2ouph7nYoxj+SoFmaMjRdANJ/PkWV2XQ+nxjHA1wJd4M0v9JcNcZgXVQ2mozTOzDs
dRoxvEG1Nq0Q7W5GRZ13PHHL1+wwlbstYu5ovTFLlOx0WbkqwNRIMtaWqJoB3Rdz0rF6vUrOwoyV
EMw5yHWQQ+ki1CRTa4YxHnNWftNj8Q0tlMFeFBjJOtFD+34vCo76lMMluWXsfENui2uwyqLZqCLu
mt/fXuI37RZs8Jnk3jwLU6hFigcFMR8i+8urXDkuNiR1B8rNSUQRjY9N2h61TCnIxQDkvjNs9woc
WhYTdQYb+xCSO2UYkPBgPZSSSz0D4anwvpgsRP2uqGWD+c4CEJB0G/OgOFqEVIRdx20/CD202tlC
tAxtsIE2rtmG8EWd1SP1Z/Z9KXQutB1DKKahOg01H4jpHR53TY3wA/U2kFzjfxVZIpgu6NVxGFg4
p0mbEE7y4FhUu6K92NmIvRzyY0QYQFEXHGYUk9PxJheTTkf4lLwCxi02A4N98q78+qw7Ig3LMDJ0
rYb4IyfBYqcYWzGt8SQ26rxxinPNgeYKObZWokR6CEPpSUVrPspQV0i8YzlqbuQCR1VzVm7n0gcd
7KmYYQkcDVZmCxkGnrmNrsAM11+YcBQ53Ehg/vEWhwpnFUjnqjpR8Us5O3v8IuEhK6pZkIKubF8m
Nr8J3RkmgWKFMPuau1ADKA10s7Ktim6PB4FD1NaJ5Q21ke4nlndujKLdeY92zoBLpk3UQ3TBMuPX
DVhW2DWDIrAuo7pc3dvURkWgObbJBh918oWwP1EUX9gXJ230Mt4whnfYlTasoM+ifQd4zmvHTaS2
aPSo6xeB4NU/3Eje5bBSly7he2hB/8UJYLo3Zb7DbreEP5hQnv1FjKDCVTLSDRCB+uBP6A1Bu5s7
+AsbzFCh+SvkYfIGXfOV+zQM5luDYu3I9h+BhyPT45ih9+UsWvD5/6Vy912TRXIIIosCAgzeZnRe
CtNKRvR/4P+oKSXNy6vaBup+0jHGwzHuhSaK/vdckMAr0qrY10TAXPEIoBsDA791ZTUkMqx4ms+S
+lD3JVt2Bb4+wvAdR5fJWCXBC32eO7dfkEBpxAMaU2oxHfJ7I1U3zO8ATFhpgr2JMw9uEA7TN7SJ
aeaGXw7Yk1CzwDBvm4yiP+F3+O3wkT8TpyrMk5VRlfan224xFqlXvzD3368bKzxlRjnD1X5R70xK
2F468fUAhxbkDiuiOfA4X5TN95R6pkcWY1gbbY63Hw9lQnNPnVFvvgf3q/3vn+8jqWoRcLXhkNUy
0vepLlClGRJMeUgeJaIPwIcIXXz+bcJOXR/j+7mA8GI5UagNnNsNNeeMOGwuSYYFkdUNRcOop7YJ
xoYFnzCLw0JY1DWChn0vVrpIqNS2L75Q9j2it3/wa54v1eJJlPyuuLxIdT2FyOhirLk8kTjWabTq
Pm29nXTkTXp2cpmuA1nK1YUPqXIAurmcm5xC7h9GRVx4kacGl6VH2+KOlrSGcgYigO41CPmJK+84
HT0yJQKn+FOalnY7oD1SFyV/EAVC1CSj8Y/dojBAayJc20Bvl4SCiyLBrFzjuzU1F9WkjvfR3Zw+
QkAvWw/GWRt2lEFhKpbYMrG+ED/SMtcvpc3XBolLPTi1rL69aNfhUluIQnkmdOcxPFVt4D8GBn0c
2v1NNq889cAz7Qrhnc3zI0q03lhetG1vmodCHQFnrUtxk/Do0XnElc6n+QW2tYw4rUQ2D+xc9zgo
jxswqdsYLoj1MocY/dYRimAlKxRSspzPYuGI4/q7zzvs6qqjwybZIg4xDoWfCNCGQ3if5RFy5xLV
sZcGohDV6pKWfCIc1ZpZ4L00loRbCfOt/xVPJjTzjKTbKPEF1CtqpWdQQKinjs8N6+hmStwCgV+Q
XbZknqcovwlEL9HwELVdNX/U4Y5Btb0iaqHP/PFw89Rk/DujAaWl+6ZLmO3B3nLzpR58x/WoEInt
q3g1Ju2iy5YYtti8CVTHI2zd9STMSaN1aECohuPWr9FPtgHoesgExIdcUP/tk9aZeUpVA+YBX1RE
ymyIgO5BdgsSaTLlC2t+5zj142IdC4Fbjd64MAcDGYba9rgOPPZ12t/im5x5NYoxhMJ6YwWpYiI/
U+KG4UW4jThXszNPHNfN4Zb8p7e6dkOpmfWKXmUALmEGE/QQOODpDJFAohzLShZQOsrsGH7ZxFRw
NQaMs7m1hT22o08NQk7Be0QPjvMYxR8+/wFwKivqflg+H6/WU1GcQ83yxdqh/cwuXC9o62TcQlpd
Ocj/qDbRyoelLs+dLX0qFONOyRrm6SANP8pvpE44bD4HwZhlnwPvr8MgGguoEu58NKxNWq7A0HaM
ejHDx2qIXTOmxjOxPyJUoPuW9TII/J3G34PBC1Usa6bp6uXTB+vD9GS22iPrd6nnfzHPc+ZHyBGz
pFmjD0xKPolILr+zhjjbyoQHXeLjy5jbHwfymtah8gNXkBE9SsnaDrsKOpV+N+P5aBonamluZnrA
RJhtx1g9mKhG5xeTO8OJmpifVseKReL/6tJrDGZcOnxroxtZzOYOuhxxVz/jukWVa4Fy9lfibiDf
nAmGc0q4LNYJ0fQaYNXavBLsywh4CLXyLujz1+3VXyHMJA13gMwvyLEHUtmrDy01SsV6WDiuFfCm
NPgy6rMbI8ejju7LoMqFqFsFB536LxYOjNFUqambAunR/3VUsYxUvTgs/Bt7SRfYs33s3A78joRV
MZAn2Th8I2hV+ooMHYcBB+b95UNK2BONdZzA+tU59YPi64dIvsFRoS4E0Qq85+LRtuOtBEELMZ/A
D5gw7Ng1s5hx7F1FKcP5uveVw4j+eHMiXDixIvD36fn1LSZjsE7+MIjgeu8AoityCgYZDMy+uyxs
/xRLctBNScpvIT6tSUK+4yKLi5ngIFPqnrWLu4KA+NX9v17UaeypvTeKTJA0HpgAW4+Mq5g4vvGC
m5geNseN6SFWhy3tR4wOY7gonPqcQ2q2TFTNHPy+OpRrK7dEZxU+pc1pu498t3OfnUzuzj89Y/Ec
nvsDk2WOLBFszdsjlzKRdc3Qgfzm2PSgK98xWmPvfpeRjAxe2Cu6/ULKJDizy770rGGSkIpdnkTx
eAArXmu1bfev2PptuclZFTGYMutkTNRs6PAS9utCf5uLB1EOI2kl2nNPUZGWuEcmmrFT+tnzJClV
lVfVLbJiIV0Vf8IOYU1oMdZKtasnvQ+/4L/YH1YV6iboWD77RF9dzS5TUwa6XsW0bvDe5ID0iLa3
oid++8WOFZG7g8MgYcO/FL7AiczcZiq+3VXbQ4uqJ/7gYQTE1G0iv/sSYhJG35mfPmzYcV5FIqXj
EXX4fkMpWhzdxGMIBE+/HxbVJ0YAoeefnV6YQgpWwzAloecObQPm6GzrAe1b9uK74Kk9uK/jg4c0
I9zV3Ulc7t1Hd0tKcIxaHByVLE8leuGlIpcIIOpVF/He1BCE2hAETHyt63jcpp4JIcBvm1zBOjVz
Mp3bD8Rxj24jQ+xhe1aYiq/0Us82oa4KzWhb/SQyWaTPnpvjyCYQ15a/HbGdjsONvs97zN1293B9
Q4Ew0p4ZDjs0/RKVbOyVRN/m38Cac13BCvQx/CSBgxR8Mn9yfAJqx1Cz2MLyOokHshxKZf6vzHxa
mQGjXul+mRA6eRXBSbfz5nyb5ech3JoHm0ly1n4S2YP0M0p6UR7vHfarirexjevgiYOCo8bKvwyJ
IsltFF7KvbRuqikf+ZoQ6HOsSucDzmwzyYkYKR/KOI85nbdjBPpxWgRpptZI/Aymipmh+ym7gLTl
0EbfgemLbwOED0OaOHVe4g3GGH/cu84Y/zAnmCIPKJhyjtz6VQKuzSWQ2qOzAlmxVe52pzdaDYtB
ES3/ne8TZeAmohDa1EItQgAPo2s5p6dJax4e5K0zC6GI3mmR8ju67PiTkyXzprr7igoOexWJenzY
upFUE41HF4GZsq/vkBr2oRdlDTZJv3ql5YeCtijJKvfXEAH1QFRNQ3zSVhi5EyJYPHsDyOq2tCYi
gBH+EyAOVYcSuCnffnRtQdWasJRakVyNR70TbShZN0pyQ7XuR+sChYbEHtEdOl+n9zdaBS5nbPm6
zZNLinyVC579xO18YN5rT+OPCzPvhxQiJR8h6gD4hLGWWsfdK8QWRiLoOwdmjDwmBbOyejgU2psG
Cw/WaqotBgqxZZCwu0x4Qu+pF5lCgZOdjvCtxxL60YkCa/x9A7pHI1DmSI0Zka5bAL4ue1dC6e+h
DtSUL/JyI56X+UdeBvP8OjaxX20tb9k95S6hYptugVmF88Mv0YJ7N6XX+p8RqXB/Nomm2wPhSVL6
vrEViMDQ2nQ5U54/pMpAG8nYGF5hnuAZVvmB6r3+X4LxUJNLFEeGx7agyibLB3s9K8tgu0s51+ai
TIS/X5sD0R12VPSEpyXHkAE1VzJrbHbEFVIKfOVljbMODzbP3my4y83HXvfE2RzPbt/V5GReBzAU
keH1Fy953v60SQh6AAVanDvxF8/vRSSCAuTz3zMRi1r+bNdrTWXtIDqddhrfPn+hmScOTmMGCz76
Qs8WLgHYZJdHjgiFOQyxqHyVyRZTxu6cY1/49QYnVmSm3EqOeWdajFrealNTLyEdsQ5/AU5+SqXO
WnfWpV7LVoUWJfuU3XJ9dr8++I6t4xjeChc7QvinfMDp/McR3azFtP1JmJvV+QEE/rZ1D8caex3b
GxchmD2Gp15wopPrTTguow+ncaM+UMt1G8eDbBX5Xmo0mtQQQA07ugEQei9ozVXfnj2BMsdb3Hbo
qsu2S9+ZZNXGvgM72eq9wkv+PyE0/O3bPJvfaEav5qC7T4++Gh82IX4euEi8Q1jJBIm34kuz9515
cX7zNeKwjTwt6orv/fVxim9bSBmxdkVTOTNDGCS+jcqJ4sFA5KFM+whcvYm4J8R4Aq6nZ4JWDEtt
MdJDRCezcpmlghu1zRRHx1G3H3CFT54tOgudigb0ybVDPItOYXeuKv/e+ATyz0YnbGqeIiRWAC0v
ypSAHOqr2D9OKh34WbeypnWDZxL4eoudekrMvXri0rk8aLB9HxI+NOucKdlBZ2v7leky5THXEDcX
6gvSdpbGKt52nBKHICii+U8Z1qIeLNS2+T4oGYcWJu2Qwpr/dRIA+YyNQeEFgaUH+lKAUhF5OmKz
MSvaV1Cn3bfqMobDeOVixxxol3CpDVURIRCbR56bN3FBY0PhrqawOKE2UuZsieJw+QzQBskADHIm
K0uXZoNSxjyGL45K0cB5iqKfz3JgUSAsHK9OvVdrh/+5xqBq1xcl6QEvEWTSMMypRhBOauelRNQj
/0MUjm7LWepC03nVlSHVGrAD4JK8mvF95QrjwFOnBYnLqfOoErSYTV74l2tyy/k+Pkn8TReXFMia
yeChJ2oxry9ruDGneMSAXeQuY8LnIt/YCd3vBQMhkVaWuZtqZqgOlXbgRuodztwTcMf8/C4WkWeR
HkB3outqpbA6Vu7LrIAVb2PAtZXD7e00peh0JyLIJ4yPQ9FeR6XueXqxMBHhMlNkowwrlvz1DqgF
rRGbbByWMHc+6sffI1WZqQVXv1Lq7Qi/OGeKJdMbf6WdxG2T3yTYDQIh7BNxn2eUFnd4ei0hJ8xJ
SZa/AwJwa/704vUaUSx6wxIYK/41we/5v8Q1wtHcgtu7LN/W28RS2S2vS+KwQGoYgqV7aogUhv7k
fkk0TwzSendFaJxFqrirGVCXuqVeJMstZCzMccS1dBb/VgBPZKANkmHniXLT3933DybGETd9hRlb
jdJFGf22QrxnDCPJHVev3eVWo8+fL5STO3usoUHwaDClOolzoG4YuTWXZbGJXaDaLvXs95E1S8Lj
3JsSrmsKiUGI8RKcXosvWxSikN9b68VCe0xOvfaRtajqCr6WFSapb1DlshhGmlxzvwjREjuT1JXx
lKtIXQjJ9Iey5bswAiYA9ejFVYYXcH9YUbolYKDb90MJZlsHdgFBpvN+iK0t+jpBEs4UY92aZcyh
SdSr4F/Zo4DpGdHmJzUNgTVksNjC4KBFLXedb+e06iQp/IOa0a/bWsKonfvfdv1Zo1ZFxgxB5fF/
5TkaSFnipEdshitLlw4kvN/TetDr8lCDRO/kCwBz56vc/Hk6eOmvUc3ISspEV9tGOTG+efaUjiRV
R5b3G5JDtfTiYlJYs1qjD21BeDLUeZTrGJLI2PC2hmvg0fm7GjN1cV5oT1jfglVXF87Q+DecYGft
vpiaCG9qDw5x/GktqDFSKhZiyu8mtyvC4k1h+sTj7uPxUt3BoGST3w8uiTXP0nchmu+ZKkxUanol
lpOljqOzvqzfnzQA8DRBy50smX3dutcMZ6wlMVFJDNkttKz10iwgpj7rO/OQtKCqXJPteDBSUtZ6
mayuI7aTut4wwF+8h6laY1nnBw+aiXpwaPecADoIY5Otj5U7HPw2Wh2dCey7RKNE39TUUj6g7uAs
j/LO2XLZ9f6OZvBp1UovPB/y9z86N+hbLCI24jjzpGu0+XZ0NQCVUN0Mr5fL1eCXkYZ2sQRXk+pe
O2HoGmdgVOlZbhUVcoJo/oSriOihhEYnYBJgMXlnIXi9nA4u773OoqBznbTLDJMAzOm/Te2cFI6B
IrW+1AXWs389Rem0lEiGoITPlKaAxFioAkS/tzpm/ac6d6kDdZ9YcTawI1cV0ntxwICtOy6Xq1EH
phnaZBCyi+gTE1IANkpE/VGmAcc+Z12lPuo5/rimI3XrbNxFvJmQeYxy50x34upsAz6B3XIT4+4T
GUZInQ/Td9eZ+bz/eqIIlYenfSs8XD7HLNK+g3uMx2ZFAE3f3M29JUiMZi0lVXtb3aCJM9/v8ddF
EN2MtSWuDeRrIAfMj6kOuAQDJn8BuTd+jRy8iTiupg8rCViIWEhfbiRU+IKObeWjArG50ncjDwTr
cOwh3jmduDB/vgl3f3hcNoha5g2TJ2J4h6A0AwN9CQVMWLs11Fpr1iomVEejJ3B4Ypdk7y3kvzQM
4xRSjTuMVBUv0yDCDvnNpYA9KBbsHjd5OLeKJgB5ffubQoQbCzeoRQtSe9dMB3YhBMCR34J3hDCf
XUr8zmXKL//Z4WFVlTgvPczyKCHr70Kk+uQT2/4xiQSnrZtxzMsj3rZ5d0X7y9TyDbu+r1XNmE0M
mew3XPFFuoASEui0gLamregr+VaabEXWn/ijM8yw1YvJ5Jl+yLw5fhBD1QCX91FlGzGMYBl4JGYm
YHLQdiPwCdpDpXgnjN/W1SK0HFzDlViadx6ultwXiAOIKw2SdwjPv+Q79CvHmflSAABaTUcC179K
WAyEbWVUQ7Mjyi6c1ra/ScGxMlFkanA12I4+Wqeb+6B0xdbmFAZ36WAQfoX9l758E5mrQLpljuUk
riZDqsg5lWyvg/RB8FJcfGLejTayywI9ZQr3GVzJV6EnAVn6szBoWQRBv1XBae8f4rzYF8GBTPwS
pKx8FK0+Lz2rij5IJCT6IErSt1aHDrmSyMbRXaAJYPapk7na0+EJS4rOB6L0HMn6kciB3OdRANRs
OPWRNYBf82TNwyk22I8YNW+6vclK7dgPT7uSM/b6IQc3r+bX8NSZoDPAx7EtJnfc2987Wg6CaHgm
X43j2mcA9/7oH5WxrKluQ/YUA3FRSVFbNCUS0smvA6DOSjVqp1atQQX4aBuV16j9ItS2Am6W//LN
jTQdCFV5tTh+8zfSko6BGdNcuLjpgF30TKSfFwFNKuBc6Y96IzILgnhpY1V+w3JUtzvoxfRCg9hZ
gmgg7fPww0kmj+/ZALD+5GUgJLTrRNqGzhLeGeXOqjmzckSly9/PE0LjIZ8V4A8W/tpKMzmrudUK
5SbxhoeRdUo4/AVrWOtWPDKQmoGwKs1J8GBg8HwgSXhMasx5djYgbHH2H0ErXmS3oU2rw1tyMGpF
SFYr3HzYZvLkyqxXw2c9laXjphFO6ugbg9YOJoxESHWfnjTb6OqEs0sfU+7TziOCSNENzRrnnmZ5
Y+ncnRDPjspBIpLlFkxnFUA10ZWBOv7Z+00lKbNg6UjP6MQSKyEMqI3kmeVMPKQnPZrMq/f8r9DE
mWg+BpORJLb1uyoQqI1Iepw8dbf9vjDOtZVYo5f0lAVBBWzM0bZsdoPtj+v3Hp3OAouQxiJYnG6I
Hh9zF14yOcHTUTJldfSFMkT31tpPc9XgZkyhVHXHDqcKMpRaOhb6AUYQyP3nn4j7/+dWUzQOulF5
dr4iVO0SVeAJQiZvlR7DudpFFzqQi0M61YZE8GRTo/DhN+zBdrwb3/8AYOuJXRgyI65BIGmm1wr5
maxBsY8nIb3AjQo/fx9hP4jkd3u05FnnL469ij16DBbSMIM9MuWSDiV/2nlpEvm3qOh37WHte5gb
1CuZjPhcqB5mCLcMBXpeO9t+4M0lKPdq+uF+BZ3CtlG/AiirDwxiB7Su4mKpNqqHZ78EU+1X9WZz
+X5VRjcRqg0Zy4vbheH8tw6u+SHpSrNPBP0Odv94ijL+VnHBU0CtN41m15C75vsHczwEqlUKppti
AfQyget2oaaGq7iF+QmNO6wVmzcmCEqOVl1n3kcQMgYPUC3TBNBXyMGb09vg9o0jwQXebhpRuv47
EoavW8ElWoP88PrLFS1VRzPq+MggSc1LJyFRUZR8sxB3JMxLg7hpWc7ylpJbXOEhjYiCACqoLO+D
NHv2FwZh/y3WBwoKPCf3TnYIoYpDhvCAruuBm/7wkbaNhH1tDWuo7VkI6bSfv9majxncqr+2CtH4
7+2pZFLFx7ZvNrcpoIvJNLadoTvkyhp1BVHjkE1npLCATsdj78X4sGsv08GfapUgL2L8HLcDH5+2
dB4DLVMI8cwCR0pldFJyBEvcHhT7EBu6rs5lZRkYGKbiPAfET2ybC+8tNhGF3LgmF0/qBFhr+Vei
IoSu56sQqXsgYKp253ZbU5jZn2uYBeKC1nWM4X9tfY1l9qLZ3iIdJ0xvKjsCPDs22zoSm2mgXw9m
rrrihz/IHC3+/OevZNC5m9/e8+VC7iYc5qfIUQyV1ZtAVzUzBWCGnk4m+V3iGc/9PBiCZgIkA6Lq
puOU/ZQQHdwboPvT6uJz7Wwh/N0+bvesHqgQZp5SviCsLfBg1xAI09Wzv8bCUwUfqY6mD7RLEja5
GSr6xyMoRmN2Z2jmKZO1XljMBW+xnRdPcDL7uvu5GSeqS69/vxnX9Rd7CJztTSyQYR8RMeISnb/s
ghtH4leB6dCriPKjk/Ydgo/mrwKEx6Eu7DD8pjIJ4EKR0Su/P/3SlFQHrIgSngATOwBrdn73VeuM
uyQbMKsBLaT83of78bqhB0LRIn9FwW+l4BjeAzqFIhJ/NAJXf6E9+faeECS2a+l8/EAo0xEsV5Mq
WSqpwpafa76rN6t+N9+F5EyrhBgAjuFvNlDtaWXOrIFCxLjakICVjJaJ4gZiEFEgOjv/pxk7TQoq
ZuWeCkkkKVX75uqJlQtobLcphIFhxIUIIjIvUh4Ip6GCm3FN5YPT9MnTnM2rR877k0+ATjI7NF5n
fLYC5BQ/yy3ZFKEOHl5FDFBkQTOG7eIZLGwsTSNQMlkx4GKVZeSvhFfoIrDhdJLb4hSN7oJBCvPJ
rl5gNPYo+YGfGRL3bcd/wOD0pJ4gn86ZQ1VxhxZ3tLlkt7etRSYvQVpquRvjqr9xlw3i2QhS14o9
SxpmVGF8Outinf3U15rid55FEL+Mg0NyOYZq/WDfDI/+d5UgrFFKaIWgVAuBzJ/6hXb/pLjqnwSv
O7ZbMgW1v30TZavWVFuiYf0E45LfUt6TrFXtshxT0Bq5VW7kjUSLrE9duPK6N1d8CGggx0Asrc+J
1XW06C3yQ575UGkoqsjYpInXDGlkmXwiIpqlykqs7Wgyw04+iKPhfxELtJeqgA0Y0cpd3WO7O8u0
4znETqVHGS+QyYDLqqPuTc4eCTGsOzuGtfdUKP5EzyQe9yiR3vGV2b5dPwDGz2tqQa22weYu5gRq
o+Iqsh7UaIJt5JgnEeEQ9nBCcVFz2CZlSQJZfRsmBOCo/BKOLDuCsVToCP2+JfXT5S1A+otWATVR
n/9A1HNYqVtIta4ZqOIfT/9qP4W55pLZD3JjPjNtl2pdWZhK7qwIrm9ScN3R6Cjj9tx5auecR/jy
pyehVCVWXoI98nGp6EjYwAAPEfZgdyQHc92CfrXxsXO4/4RKKiNEEIKD7XwOgh/74nLYoAl+b9XO
6jp+L6WE3UJQzM6ijCL+pIM2s4KW5UDXNudxmB9aNlXg76mJFIeS7uOm2cpWp0Jjs9CmgkUQEV/r
RYxGXeuh2j7wPs9QX9+7KMHm5iRuh2ZB7YhZz4SJTsINoga4KR48NIMWXSzG4M47PmiwHbC19HmZ
4bsw7IHtQTp9PdRjJmUhgkO1rkSn3vKZDD/RocNk0fsT2D17jc0dOX877gTQw3FRSx1FpCY9HVum
kJgBEckUKj74Umpoe14M0mjoLffTQyTMWQxwUC60V386Wg91Ur7jL9nxnpZUc7KbNkKbaWjaOxqw
eeVnzaGJAzRh4JCOMHDK8CBgNQvOFAAmyeUPB1R4wVZb9PMNEMiX2owcAj4ZLPozJxyUCYbIDU5C
10Pbycy5ItJKCmCOb9OAx6UA7If0ntqcjZ8p0kVBSYJV9yFpuptOS1jxxj/8A1C6/UY3ANRLFeiy
35AI6CK0bYafDuCbo22TW9LzsLEJDivQabXvgNQvT6PD9ZXPkiBa4Q4/mGIrMH1vYGCkI15wH+Je
//6b0g9gwyugayENBAkBgPN1YnidrM3l+2IUIYN/5Jzt927oGzABu6T0Vm1php1JGA9M3PDssVVZ
rIGsSCVE84wZacQbQeGAJhhIF5dgQSTGzltIClk8wM4JJWkLeYN5bylT10Y6axoKA38zBjNNcxwp
C+YMyGEHLeVN3BBzVcDyHX8+v30MJ1layuMGrNI1scquHz0XyghKEkuf/k3PjvGVpoc0TFzC5txN
RAEqFJ++MCcTUiW5FMK4yUjt8gmNsbCAaQh4YXtwuiaRlQMwnB7TsbMCvgIeVJtb7BPy5D162yc2
Bn3a10nABH3sr9ZIhZ3SKGs7kcIdGVF5EFmlxFL48aroLhf2y6OugE0/lIR2fEecqy3EGS8fEllY
EXa+0lEp9tw1y7JW/C+NRE/C/lAF5rtVlTsC+OcDfARpn4siDUMaquBbGiDuzw5FLbPnaVKZ5Fle
AEDj8DBjLvhyBeGH95xsoENwX7nRiUyXLDUGiecWuNSzFY8Ssl7mMVpPSlVRbBwRwUyWfD7PEoNm
xWBZPgRFWWH9MqmPiIWr1AZoiJy0sDygN0uahbxGQKy9jTc/8sGgCtSC5YbxIrfJ/u3GtGEdRqxh
mhUg6p5VpndoAb4iihgJIQI8ew004zt4Ams0eAJKM1D+11N3P1vX4Fs9ofuLwvtNSvE3+4qqZnKQ
BxYQjNUfrGA8+8iDeehbkieS/y/QPSOBhsio7Qk/vOodMzfVe+I5t69KIkweyFBefj/XqidFQlMp
OxTHrX8OiDRK8C0iQ7dlklzX9G3yKbVBvZMQDkG03zsJknJ71ecl/aI88LYAU0dyZHMW9VS+Qvju
N1WGFX9vtfVmj81PClB0uNDkQP4GdM+RdL/1ruD+zXqYs6dWglaoRvbcvfTpkugV0d0j1dFP4nFd
QBPm+rWewwfEfkvmSRjXBuCHAOJJT84nZtZ6BhNfGM9JEvVz2YdnAHgMJo0P1v4n2PQGsI136vec
n8CxTC0LAIQ25NQkZEB141ujbSFhHpv/dcjXI0eGdMnm5d/Ccv4HzG0jrgb4obfsgVT9R7/XH1kB
P9aNt2yIpaMMAAQPe0/Dy9FqHpUSYhCPVWrJJqhEHP3p61HGSU8ESvoohNgR7693EwfDh519AJD/
7KEFzCi7pOQ+Q+GLTvmBJL0HHHHbX41SzTTsLIcVC7LID+ROvuknE1oZJHULa6afkR70o3zRmNFK
j5zU2yttZ8AZbTMYFwYfla7XlcwjrzWR4GThaoy5S3jcbrjhC+ppkt3f8cmFfdasNzdpKL6hCWBm
5T0t7927vRtQDQpf7Be6nDFjuDNczN05R4iDG8wmzmiPBDvEpqAHYl324RiFISB9ExpgjDCr3zx0
eaNf7+q8QzBdH8kriM7OAJ7ryY8rxDRuYV8QL6kn/+CChhd4PeqsFn45rfnHpKtu/Jc2PQ2A/h6/
8iFt8E9lLo2NZ+VYm5RUty8AilKtDcqK/i8iu07jlPJYYgGSW2P+Xm7IWXcMP/pGSZIv9EaNAFWD
whWnqCM82C6oRV924sXm/mjw+mg9/ag+hbU6goHFa06yTyfBwCYn1NM2cdCRnaim6ncAbu81ZOlC
XEE+to08KRXuyYwQCgiX80q3M2NwqX9srmenPeFkuGYU4ANkQtGKbB/YJjBEKCLQgwXUounCcW9c
mZuVrWpSkcbAVMjmp75wqeBVEwcaEOpGO4D3JmcxLfVwcoRIgINkKW3y5loUMwaIVSTPPfIST7iS
yVzaEFta5q2IZcGR6/JWx2SRmCqKZK4dtJFd7Cdy9+/KH1NjweOI5zr6wyjmUM1NedWBErHYu9Tz
PC0V/BqjYD+gid7DG9Qxe61XH8rOv41hwShx5KgFIaPVc+i8OrIdxaCxw97SaIwInIAW/SDyiCPp
2FsUznsfXf+gUjO+00y+YyALcIQwf/Nzv/NWNzsXtcvkBu2M8YE6YpKkAWypZDRSLq9VrOFIYcPb
8kjWVocPUQK6Ysi17NG30YcJLM+nPXxW0lc+goSstkL29yjNIBNnV94Ty/DWIW52WNAr/DQdh44C
goC1xxVqtwcimgDiXYYTm30LHQNYtQwQ/pLE6JfdNOQVH+QfM3hE3ppwtmejKJ9/taiKL/PjKt01
PtvfHs+CAe7s3vJuXhZsRhFAY1LaqwI2WTLaGGj/11b+jrYXXAoOZXQMtZ53koDe4MN5gwXCaCLf
JAIbCUMhyQKhFx22QNxCdn7Cx5x9x2J0zgxWVJLvhP2vp9ByMZkrFsUTGktNtF5POZr3UPwtMVj7
/Ld2GdLLp4WJyzaUR/mI+HnUPMDG+lp+Mt/3SLzEo4UoEyo91SwqIMjd9/fhB308UL1jv1uhBDoX
SCYfx3TGTBYhhV0DIqd+fdeEuOsVoqmoOtYvFqUDEb7KOKD9j6wevky5R2d5w3QItwvu9GIQN8m6
Dy87Dkr4GM+nR19O/TQyrXB5S7Jl/KlxxYLWVRic5yGVuESTFO/TnIeJxM3SMfxTx/M4/IeydJjw
pUuRnDaalq8FzKceoIxWQl7KFSJddpD6yS5K+Ta2dJLJGkakvOErhk0X7G4J/tjJ7RazvDyBhIt5
ahvk4I5qlOXHp6P68AbRQUI86P/xZsCdtDiYwchxXwb6ClGSz6MeDgCpT8/oAVAFM3XkdnhvVRa2
iCXSa/VHEms3iIEt81EDe0Ou7PFHh6rw/cm4KfyAjb/XyfEooT8+5WoGP6yerYm/pSaxIJ74WUk5
SB6EZz6iSbHosVDtlNUZ5g3D4rWaIDYuCOwTG6rLXqqBjVS/f8oeQ4YLyna8TDdZi6w1phpQZems
qgjw/45K06dBkB0MSOBWz6UCmFAZM6hHB1o/xvBELKSmmjxQtso81FcLIdMkzXJZ1zrHqSRbbkLB
sJyMBgHVA6dbDn05HT96GhcqlTWjOKnHwwpLUjR8Xpo/M9UH6YnKYBZhx3mq9DsIautt79HZNKvI
PMDh+eEf08iRgdbaAoTdjEcw4d1nYt/ZCadF+U2MvlAAx80X90CywBOmbkfDu4rDoLlwFI/d2e1s
bgO3msR9+lCqMsDdPa+KBqKMSjSCnS+KdSQ0UZY8+6ERKCZrVDdQM6MW0EOzKUDd7h3SUafxMIwJ
Y6w/adA3+sOWOenJprr30hhseKj2ms/6rHHrsAywUvMqhEFyrnyPzY7ahW8YrVf/KxhRHaFeAHMX
XhG2k9IgdcezU2CWmeP/de9ZIlVAAbDBkkDGYWsHONGuOtrM5SRHiiQ5HMu26+ykNbSVpZlkp2z/
OBVbQIJnMM8z9DtmTRl3tv8A+QYLJnciGf/WXVIBk8PHdsnrp2vUlJ3pMDV0OWTYWVoWLT6DUHFM
C6uueM737ZrFyWu2PCjrSAh0FJnu4UQat9DoDSz0U55SpsCfkFR4yNO+amL0mEGF1XgDpcEI1XFK
Pe8gck37YcjgMQKWLLQWvI9Y+gaODNgyEhpFTjo39XYhkaZTg68nUT/qmt9PCMYkmlCR7vKkwdCH
aOAse1taHiGcKw3cceav+IAbgaIfnKgJta1OsskGp7If+2D/oTndFxjyxopCzHdJXI2bK2xAowJQ
wyK1k6LxzSchdqVCAhQ3Uph0GMoQ4/eJyaiWfR5x6W9Fj4JPopuYG1YlUKD7HL4Duv7YYgwdns4H
ukuTL2KDAjtlyYcs1isi66pDD/z/nc2IwL4NQLt6xk9WWIu1giH83XntGXxorsZZdMdH+KXyQ3uN
Jq7AoeaQbzCzF+Pt5oKDoaDhaDlSgDFKK7csBtmndwmoLG3tfCftwDvo98HChVEDYCencwkIYvpP
JXDydpVe6TYEILd7Ec32t7NZ62n2/ykPyNLGphKfzRBeQiD2l0FzhcdY9TxGYdAJxRDhyIFadkNm
mI2ucKPTHtHZ0AFKwikDS1UHlfg1Hmyg8gmvSn7ZQydqYvGCoIzG8wp42dGjJgz/lGAQ3Sd+U62n
/ObYUArRvmO7HUavDkwPiwF9bhaLF8vHUMtgedlUmv2g3K4gQ1YZyJGMOAq+waGGa3tHIV0lE4b+
BXYKfwgUO2h4ftZv1Y55NOEFILW616FeYMAy0Zt33IGv3AOEvT/EHtGYfJqEbMdswyFgVp7IGks0
LlL5pYNPiMyjFdQ9Lu1x4eAZcPGR/R9CqgxMorWewXRCWOHsAtuoM6J+gfPgpG8U6NB38iTWAOeT
BYxZ5pduYvgzNaIu3efZhLK5JEHz6wOEoJgulqhinWa3ZUqg/kWnlkl53NOY+Ii+ojWU1Yt9LyaD
uVuWhfHn1xKEY5GCLw0RuUIm6h0RtQwh0VxSG6z3OliYK0WU5DpMIUumXcnMx64Fw/aD0a/HiTsF
f18b8jZNbx7gM0Dm5Bu9S0391kmeXkTjhQIddCjNSHWKKrO9ZeCQOjO9ofXGA4x6yQK5/1JSc6NO
5VAoVePC0ls2M27l2wws6L5w4b4OXKjm08ihyk+JNLszU35sOOgoMhYILcz5fZWojuP8mfcCp4rM
lZLqQBUlhXxLpyicegZZKPiQ7c2mqqZuNNRktymxLnsd7KB5vQWhjpYvho8bHmh3sOsWUv59v5dP
K4IVN0452sSr34i285g8rL+dXS4aQ3tbDkbzGdPdW9UYq/ODY5IcOoWG80O8rhVpySUP0pOiyH4I
8vFZpwf8rnNTi3HOWXGPN7Qyr2azO+ZSjQd5tOwkFLxaWCTDk6UL5amoWtTinlpku00+qPOy9lOX
989T+zzfGgpsp4vlJVK33GrbtKmrLGapiTnSx895Y1TyGcrZv26BZDHeuA0AwQ2xgL36XOQA/hdt
20sWCcQsp9dMUznNZpi5KVjQoFzPCWeu1tzT3OmTLVwjspsmv+kY4hLVmA0OgrYlW43NrTHBitdY
qtt/c5bXgD4Zt3BKJtQV9/EuGBG6vktp9v7hHzZLDRO/K0B+MFO6dIe52aQ2LaEqVIZ2codir38O
zAniq2KllVjZkqHRu7Np2RQlV5vNva+ytAJHCFVE3/LJGVresPa3papX9Bp/gtcl6nzydNSXCfcs
RE9DDK5VhXxxrC7eAqUOUdE+S60O3BCWlotKbU+i9zCZ+1e63dBO0qItbmEBvP6k0h/vp15Jrl/6
17+s5qq6tKi3DWViQEFOBlq5avFEOheGFYtIHR/iDdXQZTGlSX37cB6vDcP9WncD2HEOErsNph+q
hFHiRGMobkoKIxg2gGQ/lx6X+ExAylLsCp8JDwH06+2Q2YNUutijP0jrWqyGzDxVGMLDOli0v1Gm
uAo6rcCCaooYGwikagKdtlNVZ0FPRdW7xr+tm1MXd9g7+SlutXUGR71v+tEzZpQshZ7Bsnli8cNS
1R2dBC/4BK2Lx5H6iZHCt3lobaKkm7AobmJFTroURq2D2fi/ONWcUKdntEf17TnJ6to5FOO1uPrl
pVmLuQ5d0vPWHU/zg53L4DyIfzJUcLRBW0X+FUgxugwPj75l9a4LUSjmGsVwb3kIa6Ix+NRMzCDb
JZxUhJNzq0zaK6hRmlAA4DglrUAylFPeTXlnl197SUrldoYzxX3bK22OSXHcBoOHs/X/knyQ01XZ
INjnIX3tREFGYfdLMbjMs2hxc4bN0iE7YKagNE+/wXmmWjWZTlAs4YDBdZMqIhRlPQqDkukag4L2
tXjc8BN9p7GD1qV4UKjOlDqIT0lKhhOwe1kVb8oEaYBR7pmFiqCEfPTToZBEBuwFoliqgRAm/MM3
E9pr2TSn3oCBinBPIEI2bxEc34f32O8s47pNBv5A88svOaDkWE+RhaP9KEwk1tG1daWJFEnCGPUo
YnfU8Vqlq6RI7wvytp747q8xzDBL3tk2iisz0ZCkTZ0JOYSkKeQN9pAPfS78EFN6NnF1pdN3lvxR
5cvRb+8knsoOjiaGirIMuVKZzMyjI/Frzd/J6+z9nGjyMuzdiQa7I/9APK+Q6itrTX+VKyzHDm25
M/kZ06u1LO5OM9yGqkCmIMkXF47VBPxa7Jlb/kiDq00zXRw1ozzYEn7jaH64yVQBokcxUe6HYlPS
91rCeeWzuc395T+0znpE6cevogGWTAuIdizx2hiGZW01qk8+zYFaTgMqRib2ZZBvBRLpM5bXvE3l
UVoa04pmfryrbL/8ZKX/MHzZ+Bd+iaUfmOjBgkwI2tMJhQzA66TVGbI7IsgqeLVeHURP9cK/+QPq
yr+DfWKK2iU2LK1Cfg1zdD3gFVCkaRfV67o37Ewrd8z8o8IJor1sUW1bez4i5zHu4SWMIvpZSr1O
dZay6XaCTYKQH4MD18nqLpu1KiVwjH8SnhK4TP/vl8BjGosg+8x02qINu19zGX+xuqPb5yUX7n1U
zE6FofYW3OzrLE2P3I8GiMUuhLQhzvKvHPPAFp+w3ESvZyTcoOTmqL5asUv6zZvBmTh3d+65ZpBo
k3Zp3gS//XtAnXzVwpju7+6VGs6vN9y8qkV6VcdDxJJtr3sCe37bpEzc29mdroSV2cKBwImuvqVG
Od4alxS0vASefiS+56n4B8F2x0LmogzmodFDiFByLNtRrixmNYz3QGlWaJm1pZOLtdx/41bxJsOZ
/e9M93n00GAl1c5EDi/YHlDqReI/cs57OGvld3GGiZUFQvluvOnj/NWnAFfYfquoUm7XT2v23IWG
HYTpgIMaLIeXP1D/lpu8wvV9j21DbDjt7DYipFTbqPjpWcq0y45pdKDh64agpLJx8g8V/ow3CuA8
glhAjT7xmtESEFUj77V1rrKLhNB3Lg4gGb3P03XqrYluO3jVF29l55mYsYPilcxG1q3zlBA7ApI4
iIJ+guD3WHljZB5dEg/RXixr+LCD/EGz3tCaj9+O3c7uRjr82AZk0EueuJpkiNO4t5TMmgyLPdM+
1C9IddInU/9mnhxatbbhEts81xlCcZZsJn/WgLBK2SKopZ+YskE9Lncij+BXynkiDk7uyrGg4yI5
LwxMIKfldYXjE7znLujuSh8kSDJq7fQp1Nq5tx+OzS4ah1SGO7sWOkqedgeCcFmkPn7PNvsYEQB2
bRE7u3mcp37n+MlbUm0LCGPIWsZIwE83uUnnCsvEotOSCkvcTDnKOwiWsXSTYZAs96PotSW+v2+z
xyToEab2xgiikfzlSQncZ3YqJRljQvkKXR/bqUFQAZUx42O28o0s6abPk7xT0WV5MD8eOo0wuqWv
vg/y6xFRBZf63poqox54jovQrxz7jXeOknjBA2tTAElI3bDV28rTB5FnVmT23RKSMkyXRehPFy4Y
PdDWrthOQMzw7P6zlrGAUPZGOGPvNKCPL1vskowbEauQPJVMPwd5k9EDWNVb3hOhc2CvYR1Sguso
mc0qOOPk9ZCDIVq9WSRxk+XOdiKtDm2YpitW3KKGM0pASpNEIGyxcuIEsPZ7/B6XOT8fZhFxU1q2
kQn+7E8QyARlUwRmMSpN52VbHqvVwBP0STsgq31T5hEyfZoHaryYVT267KnhtuFjU8pwwBsVemLN
huaBq6kvXfWZaj5qLPqKzTKoUiA55AtljLmS1jR8bpZh69WuHtqsiIWVMT0wr0OLIj5i9VqWhD87
ATJeqBHPZLa4O3svzfsjikMavtLsje3e7EK0pKqyuCoSEBUm1ZumkqM1UQUYhN6vyynU59Tr9UDt
Ll9PQ/Le/eFwheL98QKQXcrTaNqwxlZW/C0S8ChIIZkI2+E/JfU4XKphWUVGthWUma/iJ54DnRF1
QrP9oiV33Tu/bvv6Cnf38zfw98LPEAkXDQKE6JqSlCch3JdiLhiYMMILmNjyFgCcEwBafg8h0zco
vA7nBZNn8AddKf9Uoydt96pwdP27z9NN8/ZAE0GlirLvh+pDKZr2GEBOE7huBWVwaIM7wJvg6xeG
v/ZzNefmPivHS1Vd5xEKPePIBdmvjHOCq9zxkcKKRbVxVpQzK2aTnKuAYoIPmjIDAUvbMmYS+hCw
goA/NSj8mplL8r7ySLqfavnlj7LAga4ScvRepZa6al5t0eE0t5MW2j2X38biU84Y0vSkpHqUKWKj
Bz7ASjnoBYGlIVpc9N6yefXXVCWlnRMl7kVKb0B/oUJfcK2WrL8Ux0QzS/rSV9JMEmlgU9sazNej
sdyXQdR7VogTKnQikRwDKNKw3MsS0C7v4f5AfZWiYTNFmtOEFMwPmAeZy6UUu46frKkF2/ok7kFn
3rDe6mVig6mi/88Jp1JYj7xYmaFQpNTSZB8+shiIP5hlLhAvLANcp6N7b7Q9rdyDlkX2V9zIRY13
McXDVv2Wz+37h9zvVaFt2lxCS0vueuhYs+BM0sct6PDthb40EJL4QP9JI1gDnIW36rVU0PjS/iNG
6bY01/hqzClZf+8ejBoPYyIL/2TaJpbwgF92ach6XDNXUU+GCUP7JZhwceclnfKdf2TwGsQI414S
R6n9N00mDY9aJAly78nZbTh80EKdH0F6FKmhA9Rlq/WAnqnkAggH7h91gh973SdxgPrT58/I/0VZ
DzhTc0LZEM9rKZxu3FfJ7IBDMfWw9jud9UfWQp+n+0hrDAs7wy8L2ilLT4RLqqmcU9wmP+lNbEYB
mVSIIWAu4NL4fo598EuuTRIEk8/L9RAfVHoEunBpJmOOSpelfZXL+udSLde6k60e00soYJxY+WEw
BN0QVKz1UBLZIGm0vR7weNZDuJgSTvQ+EiEYmY8dFioQw9htf1wYxQ79G1hrBgEl8RvCcs3hcYcx
okAkobjUHdwplZWZCMhL0zdvorKP4HrD7og+ZcK7ynF4hiIYPfLdYTWRyLPkN5gIO9z8rhtAlnM3
jm2PU4PcLVPQBIHVymXh1NO42QJJR8MwB5ARxKg3JCdQJ8P6V+Vz9/M6jXztLq5rm5ivj8TSPc6M
c/QqMLYFrhttVuHfjiMgTky3XZrcEpptFhM1SoZFyZqNq9Imo1zqPv21C4Ymy+HABXXulvKRvovp
C455g+6cXlxcyy/7REsJZJ08JmGixgUPOz3aXbmzmAZCH57aMUDDHOZgvPJ+uUQ+mbrEEyTRZMYD
E7Jg9UfGOUXrrF9qILdVOyp6TExETUF1KR7sCzUwCStSqQ/anjTCPILvHQAcM4rWJxUdoKm3EF0f
4f1/BlWzyhtGE6eCYnEWDOjFxRnN2OaqOKs9BX/MIHk+BcVYbu90kSOFlmeqkl6pOKzgV5bP8Vol
pZsMnbbzumrhV3fLA/UwFlfMNZCxS8nexI9FydUkUxN0vLEWqEDYzxOFoAbsprNeGkbc2aapifkJ
W5VX3G0NI7eD5uo94rtLovu9f2gmVTq/pEg7Bi6qWXlpxutTbE/16/6VTf41vN8nfZ+MXdqy9BTP
1SjDNUJSCCAv2Qh8ZCyxIiarcKrKTUtflGuFyWuleCED3l/hTkD2dkGZvCoMF6xnD5IqLr6EnYl8
TzlMJxmXfGV8VuI5Bd6eLIx1QzRp/DXf43dcyBh9wqRzgJdw7PusxFzsEF04dIFvcWMKfBaQKvg5
D49+xJLXFd5STXOBRSyMoexY9VaNuONVmw1GkI9XZ/woKIZnav8DOlN5DGwlQxx6G2mM83/EZPdm
K/lTEVAsZ7Jkx3ipLhEnFntQ7+OYvM6c23YwBNJFrLSNSa3GCFnD3+9nlLpHm8iAb22FmnvrviQD
dFB526aN2KzmpnpopiZMFQZZDREN2V8G9MG2qiUpK3S1mtVXM2OFgABdLUf8xI5YANNHf02n+zhs
s1ukNVzLbUqHhapl5rAQdxntDqkwXlXqh6lu08i9Jmv+OgsHPf9WWze9HhW494stQhiqqYrY37t2
d3VK9qIZVEBU5TK/da6wSVlhlu3Pgn58bQltbXYSXzCbJRVL0LkOOt6G0qjZUQJIXxEHgTvMoiqR
6fh1FifONnzqvyNcU5LCt6pxusNU9wmz5enDtgABqW6ql0gEYGd+AsHLwj5FxNRGN7z/huau7Ucj
9ieQqnz/iJWkhUT5TnUqbDuXvQ4ET+RgdNCGtWMbSwdCQlfQfvnYhIiRPeGbp6XWtNCHOHkiQwvF
57AmmwGkmJ7s7eRYdNW5MKuJIm8HUl1atrrJBxqrZmyRqrR7Kt1IeWFZ1ggXS5ncOqKgonjrCRUx
Qq1go5KnKpu3VQjs8lZ3RtzjnKk15b/bnQUn6pKIgtY6RKyYnyH01AORHaeP1W5W5nNwEeg56RTg
K+AGwnEjT1SR4OZ6rVKXETC1JgNI0EnYL1sy59n7UOl2nRVWVZnLevvgDptKzAM5YSbsRDNb3Q7/
jQgZcrmD1gYdT9NiptTDr+XQOOZ9AozYqUz+uU3fcHQYLSEJn+mAMgd9KOENCVRYZ9n+c5iNN19C
eBetPIN5364FidLtAPgN21Qog/45f19ISJu2jdeWirRXkSvND+0a/mDyb2R1epmYK7xYN2L2Oh56
qjFEwzKFU/FhVdk4dWQeHdiz/ZQjXUtBaYt6C0jqNDaKzSTV5XZV9PfGfZf7FzqgWckAtnJOlUGv
UeytuwZtF1tK1fOH1SM+49HMcBgKQ1mOD910ldXKixhoZFw/x+H9jR42mMYHDzRolFuAYQO9/i99
4Ia7RQMSvOARCKzSIYaL0dcAj+sPjpgZx3pxx1NPjqs610o4Vw8mHBvF1zbV9eSuk5CPhrO+ZSSf
YyT8CM8SRW38lvFbSCZLcJNq6l46e6GRDGANdVlZv99XWVYcyP1sW173r1ZRoCRJ8h/EbhGWxKQP
QeW9XBy+ClSfgFz9rw8rNJV/XTm3lklYt3z6EpshrvZy/E4IkmhWmMhHUbsX4J8J2wNKzmnZbqQm
qeYCuERxbJ4CGRrl3LXKOC+1hFnS/b5o4JWLlhEesENlNLZxyTk2K/55yr5+EpWeYFJCFX9wmKAD
oVrzToLqMkX6O76fHoIZJYqUHdw5w0a/BtU7aiVtgfYugfg1nkKw6eYxVvrWSryVbJ7U90wK8a9O
G0g2DX21AvrKlvyZpHO97TRz9NyBT5doweGBCZE3BLmUC0yhYpL6N2xkg2U2tnj2vmNK8OmK4vRA
zGn3o1flstaB+sow1Yl40k1+TUgVQrQuN6SDLwkPGrEdSdyFEwC+TnWpdN2RHwX9NzkiS7sVOjuD
cDu9ggjKOsCfbGs+/eWxHU+njExPzfYTDrK86cE4T95YO5IKlLzs9LMhAFIvO/12ZRkPcOZ7WTQM
Hd4FFAW+cXMGW7KFZUtfUuX5Q2EGpDnfFSm7KK7Ns7F7OXJ2iia98oU57wwqZa40SS+o9tlcxerr
RXmOVXSPC1uOv7Xrxk2ne3/RyHa0icF13rDHbkZiHcu1NUgU//qhnQww4lCFNNRIXXgfW1C9Hya+
ipWu8k9EEDjq+XBVuigTh9BoRhKtj3eC3gEWUn/oDyHZaLnZ9HFBKbVrwgvotDRONwd/G7/Giklc
LfvrBATClZAr8rdHQdMcql+TvSnBtXasQ4z7URbBpC+Wb13hI5RI7aM4jwavXt42nXX5g2WC+Rrn
BGo191G71kXY97ftwWeeH6eba9liPvCLayD2SKKDbfHKQMjOux1AmYp2rAQF5n0+2N4nqC9LRHTI
aDbgPAD4z0ZIKJprkLhCnSKihUZZujUtMc92uvEKNzGemzFD/OSKpz9UwgRQ83D01UHZC7BKjTXC
aJOxWSjOGq9PgKvWCwrg+P+btLfMF1SZwkiQS2sFO8V18mC7rZ538DckerX1ycaufZR8eN/za1ad
lOQfg5bkNmWKzj/0Tr7hPyx+PX0C3a/9HoTB6xb7JD7Y7maIC2Lg6a8XCsnb7279h3l+zgIAa9lw
lym3QHTzegzcdrdc3K5T5aVfyA1l2Y0lVKU/D79GcWioqhBWkyD8O3yuZb5OqpIiPoZ5JGqD3pqx
NPfRKfVOQuUnaE4WPsKUbR79XOd3iuktC6dH1f5drCwMiDyiB2QBIV+mSo1VpPJix09g5EDvPnQC
xkwGH7+XSCramK+SvNRsVJbCBBdbeUd/AbsAbXfsEeOb/1Zl3hR01pOTvdezZYrmVQs3o5iB5Wq3
583Q3y4Eg0rVqZSEzqR5wdMiHsarA86dQTbIfzM+MLp+pGVsm6qAKu/4IOqQWk6jrjLYFbwAP0/G
WCyeXupFUCIhaqKyVFM7pZFBlE2E9eC/MPfLAPVDJFffIPwctcVNh5EkXjOFd8LXHWuX65PKvz/Z
GYVwQdIYZp8o/vNon4gzVhC3mIRqUu8+MLNHOLuh7umEyyDOaTvuTMuN7STv6vJelCBWd5gOXDc+
pODHdOE7uIia4LM+fnFvlGViaiT0fKddA8tGnkURqkq8vkwJr/42CkzQHpAX2wAoQbty+w0TZ/Iy
+xDkOKBG/ntLNXps/zKpVLck7MXoB1n0FqkAyaEJ2mFExGSU31tDGPOBY/Mjcm+lAwA5N3nL8djB
7eywUIhYuswzT8IAYGXUjRf/LHKwVlgxOh6Tpmka0o94Tpirrr/wlYxDdCnOddikso87A1Onehdu
KBSe9sR77PzXYRpXKWwWeHysVbQywQOJIn7jqUnZh3wqEm2a8TTHx59RRn9plJD8YEjXOUAHqZ4M
OqG9Ct1SaJlYhC2ih35Ad3cgVLF1WoRNWuv5XKyLMgK6bVs1oBDfPVHkKKcUNU46zAFmlEL2V883
AxAx69qJ9G6f+DYPF/PoyHdHIPOnRpXv2BnKZLpuyUeQT4//m/jog+dkXwkDG8cHvP6cacpgeyX/
uVUcli7ypj9WJnwqDwJUEW7g2Q604kf9D1t7NCYU4cTCoPVpItVVXLrKq5ih1jULNG2nHWWyJLp5
7h0z5jXd48MeRU6aINkROYWGklNT3GP8xPGgZurAe5trfArL7vAOUVYoq0B+fS40D1LK3LNrtWSS
GyUeecXgvvxc9ZOTJGfzHQozqUO/dnDd+6+WPLFQMNhBhoACX52eggxOe4OiWZshgz93Iu5HMugG
37fqPSDosmcWmBtQbvdupUB1bFF34zIRnFTj4EhuGXPFzE18h7lRld1QUGKwIhJyTHJ3WYLC24RF
bzb73fzlcik7faucQH7Tez+hiujj6R+VGCmQvTApeZZn9zoRZlXcEIn58JwOouUr5ltOqe60zxur
4xGZkBdOuVjD7hHv/+aamOcKniQFW/MOhz+jxUgeP9t6VhurjLQoHLm3tF2xMzRKl9NkkGAFnj9a
71HUjBCIlCFSJPHIXaKm5l3FKYDGdL1PNCkaJQ23KwguLJelQcslgsmfENnLyL6DmT6IdvE4K01o
IcoKCbrfnRCEIqK/g29YiBjlmictniUCuQ9kyN4wm/tCPw+/Jmkl0x1EZVhntblQqF65X4Orm7W9
3psqXOmlwMAuzYnRO6oYeaDH/dj5F6JJPfkkeI+IZJt9joRoB29tyIJnyj3lzspvfYWq93sL1tHl
kGCJfjBAfXgp75oItLgtWbTDX3sio+N0DD6VkNPWLdwer1gRP9mnqm+AWNresllPB2WLgTDabPtL
xLJ3XtUOVNH0H+ubge9Np9iWQU5heeMQvgd3yZlzJTXc63RB8wXUImXmZ45F+ITR93TTFLmEE68u
E+BPQ5MuFLm4IuHXt2S51lmJ58GylCSkIRYZ6y5UpwVI6buM/wQg4yV1n7czP6Fxjjz65/gxrdTB
I+aOohY/ajYe/9fy3ZvQy6H/m4rJwDAiuua3oMLAQJTDucm5jbaUGGmvxRHU4sQRFC3K86pK1jUR
SE4paJQqkKVgtkxEycDshOzWZjHeZ4QuvdQZgHx43t4Zt9oAdCEyXH30BXcVZ/8r/654CVZHQfs0
rXUGorfyOa3vVqbF3d+GjEPoMw8IeLYF8Jiu8aNTmKrdJEcMzaDyLulm0rfNzOGPcpA3zUXpvcWv
WMU3xeRCOFEf8QJF2oBi4wpl4AFNu8MMjQBV6vNf7EZUz/NT18vHJdcq2+x7lsA4XI5yUA+NAXOH
dUWCk8LbxxgoFXsO/PnFcparnnEcBa48qNq4mCZPWX9oDfDvo+qdwM3AFykTFA1fJok9iwjitkWo
zb3eB9RMyTcws3wmWEGJaFLAU+I03bnZ6LoPmABXjqWH+T3yIGTez+FOM0/10VGlB1qU332gm8a0
9nJ6l3j877EN6j9nxCVHV3AM8/HmDQCCIdAMZg9sgZyiB497lyL/KerVJaOi1frHjxWiRx3Q3vHr
OczYz8wntKwpU1ZVsuSCtcbjNvKj5iADkK8hR5BEFhdrjpq0yrA8oQNUzVZ8tei1gjpxQmbIjMT3
8nFETqJVq6HZ3lbVYvnyPZjjwMR0qZR3j4wrDQM1hCI2AWR+EY0RqE0m+8SlHrolwt5WqRzbKjGV
HPkcboAvp5op+Rt3wvIopqq0rNY6O00Txq+l5Mekhqf9ofVVtX9joA/lUj7/FhNqXFK7uo8sT+GV
D7K2m+pHandTn5Y2fF3Zr4kQbkSlUcDbw6CsHyNEMzJ1HuuTWmw3QIL4k2MTZTK+ExGiAtV3Vs4k
OuvMDVRkgHu/7i02tX2jkq7tcs7oPJFaOZKHvAbZ7MMGoQIR6QGsL9BCAKm+DQEdiPl1I0v2x3uL
8Qy/zTMbmISVU+BX0/ic7LX2IAewFRQEckGyPrVqTRgFuwFkB1WfyIvOYT4qa8IajHpUfJscsky0
sMTRcfKE4SfFj3n96b1oPzevMnnUTBNrWYbp/a9L5AQ1kjOk20pk1PqtwC4LsxMzty2fiyO3/m+K
UUah6JcLhcI50Pgcq6Y+3gZJs/1O4wTkP3ocsCI/35bCnsGo7wx++CU/K0NQn4vwqLP1KwiIdSqO
KqfRAWF/Aqj/KXTizOe5ao8HYGm9UwYB5cDSH63n1+lpLC8MT28br3yw3mkDk0hhF+KnrlX3enVS
BBGBW/JJ7VvS1pVblzWwFPOP2NqSl7WPP60ux8eTqiEUfqe4QJJv+ZPy07yZRgE0uEQl+JMgBt0z
kF3/HgdwCVX8BluT3+/CzPhraByfPwHrqF7qnozjQVvabm6qVWpW2TKCOxmOIDHvTGmaq6sXA+5u
M3N+38tD+Hh0tE7BlSJuJsynUjK6n6s47LdsIoN/RlRMwDVrr7ybCkDoZbz2F4goD1RZtoZjA5dN
8vlaZVRwHFy2GP7ZUuhJhAxGa5juiVJNU2etBULsPXeavtMQhf49z+oWI519XnBKa+QWwrs7dRh3
qPsI6KTevpHiaq0U3zMM0pfIJ/44fbwMdPb7qyCKH8vZKhoqBw5O44FF1pMJ9HjuLor3+Pcc1QJm
I9f9OzxpfPfO3TLIJpeTFLF/Pwz4bmjp76pgwRSWcgILLlEu7RFgPja0p4RXyT0QXfU0eq0FOult
4Se3vrM2HzpWdYP/TAJVQBZZfRDCMmCCnLLBA8E+tdayHn2vHV7QPY+iovMSsaWULHROSTjvO3to
rpA9YZRGkFbL/kzMtjW3iuLLm0ryA4RstOjjlldQlnntRvvaSRuka40HGpmaFqg+NC0E0zKHW+ej
tylyuf7irHzder25ROaNFILZQOGg7YhegLN880CLllKShHc60018H7p1RKr5cwC3zqSDj8Uhl8Zn
rcvqsW2CsE3MXYuhFS/LGDkQLD9/Shebg+j/Jxmxbo6QG0vKZKJuujEhqRJVT0FsBjinKz5AuCDD
G7lQa5bd7r3vMrt3CymkE1IqyK0r9rbIeXey6w3ear6QbQoDve1cug177lbx0yNN5Z4qtWjnc0Qc
hEgwrmQzglVUZaxp0xPTL4dZ3ln+7meaMpkVD/izNLDmGN6SbirEpLziRPCQD7JVtS+zdqRhvwLj
5U+rci13jZdnet5+9y3t9WoE0FBXQtdU+KAGWCsMwgKy9t6YCbRE65XPsHyH/spiS0kB1q5gcm/3
jMXfaLoHbOTeeQ4XoBTNPdhkdInaxT++pbMaAWZhZyF7ognFqbTvnLUwkm+LwkY9+uaq/uJTeKoG
wqGSWYco/0F2+IiOsCTIDuNRpLd/nxFILNX9o4dZHCpR2r/rUnVnCE6SOlkX8LdFMbSO17Rd88dc
bTvx9Hr9CWgLalCUBEp1RPc4EnlzXZLMHz1ylcSSfpmTvpxQ1hu14OBG/ozfd6T+PnxnZmAEDcOy
HIAl6h9yJbJ8enhNuKfuYjZq4wxfswsG1n0HA0d6WLJNdtxbkcD6QEkLFkmf8DqZsgMCwJPQThtQ
P0G5SHAdaczyMZa/NQUFW0pFaOO1zgCMmel0VaoFsH4DuLYPODnQYu+uTCc3PpKi1H62IS0tuCxS
d+nBvce4+CtpXbuEUX3EecYqGI9Su+8wW50fRHCVrhM9BjTe/cHgFBB0j2iDxAto0UrlcYaD+GMl
yCjfR+t/XN/PgrHlsQL0FsSwrO8fWA7TdkZrNJ+PCT9/lH8aU0Zv1nBMjG9BZDm5xS7oCj4mMfnE
vxq1tSOd84nLQi5LDcuNfWV9zBlHEynKaAzciQTU+COhNa+PcLydw1Iya+4u7SNR8jsg1FKWLdI8
dTvIYOfNoes+1yeS/6G/XkmHiWxag3QrSeXs77OFyvRd9Xp6sfYYSO7QU2mkbAnOOdx/EYQ9JDwk
1k7ZlKV47fIR+mFWrMldLjpSbrUbEgbPW8h3iRsURgl/rRdkThsaTFAI8Gacl/82ak4ZIIj2gncA
sWRxtqhmTXWPPAN5dvN3IhyTGU2AuJ7sayOATufoUlc6UUFrfzuprB3ZRZiLRoID9u7vR4qaB+jq
kpFTvSTvxJmOXNYj+Pcx42P98yrWSgWvTV+pTp1yg+3koQUrSSj0Vf0bdYYjyEw1cGJQtKZxbnW7
tmIhDtTbj2Bv6/ve5kVg/CEzc702KQjyYehrBKN5ksxvKW0n6LdorflD+xmyIcJwKQuJ+/EzCYpC
Jox7dov2e0mJKD3RKOCjmfKyLrZkB0gxK26I0rg3GKXbH0tTWMWQbY0GB2/FZWTUcNEkb2KeoXy9
Dm7dTd7L8qpzSsBz0t2rW1dMYWc9gD6wW3xWQvh2pr5GFq35HRvE0F4hLTyi8cNUOmC8A49URnsB
leT6MK+z5AUhAee1ClCLU4+aqOtwf5nEG9wYnVHyyI9CXzAZ+5vMOcvNzle/1TyqhbffBfyr9mFp
W3JkBOSyAzUM1xTpDhbRqg3Dlq49QMzCGErqxL1+7I48rwxSDzCGP5M/Q+vcBic39Xog308tEReU
+FiWiJumYDqK2TbLTM3DBCSvHpFC20hkldfsmnV6ULBhg9m0costB3GXx2Vkv6UC6rGSZ4GHyT2z
U2Q2VFATd1PrMboi7NIdVLSGFk4aL8BAyWKYtpWPQ3+YIDiqUN6cQEl8G0vpI0/vGDp7Zslk8+F+
RFHcTYqALUL+on3pNC9kLR3xiTtIohyMBzl8yp2Z667PdhSNFVd9Bzk+VdGsCTlN5A1CYkkGitBq
QC4DtinbLMRcuHyYK0MFHz2AT+xRwuJzyvTdT/DLeFvylosu0jrYaOLRMnwkb8zFNrRmhgxHXqGv
7NIpndst6Tca3wWfGXdQXGhtyJzJs3+DH8sx0362jQ46szNq1HBCz9taX3vYWM8U3bUsnA6qIW6c
mSPAxhHKbY13ATG/ouBLHYhwDG783ZzOD6TTo80/jcwY1l/mAPXKUhazUa9mo10Ayh85CLmDVNm7
9l91KgN0nHaY8a66vC3iOu5hN3gHO5umSS7cN/JlQYsKs3O8ejRlcM10EqRFlEsxIy6CIr2/jNmG
gegtg9gDAGnva4B5F4aceKbrlt/hV7zEbHG41GjkolRMmRJkGH9sGEolzQsrNRWSkW/sADN77p2b
5qxBTgVkps6i6C+zWUxFLuIq4RZcjwxnk1T9OLYaRl6Sajlt4hALDQSBqGlOuhdd0v4DUE2yeTwS
qN8VhWxJ9OtNUjIce3Jx+iSz34N2dMZyLHPwRc3MFAj/ya9MXy+cLO8zfY3SiI2TbV3EbAxn6b+u
W5nV++CDgkaOMHfddjzLWoOGXHRrwPiEW3PIEbS/m1REoG1P+xo1qDe1d6u6Io6pqSkBxawKyDhJ
hZSaToIFlgG+80PVKupbfIqijnM3uvQztGpdoPQEyF6cR6pNsIN55m6H3QdffpwQAa5lfnQOcCch
Un9j4nmorf5oR9gj2CDVqrrV8XVjGPrhrZV5NkDV+GoOHnzhx2TVdyWp49fHHVhiaU+Sc7zN5Lej
WTG8exWfr+XFhy+cI1Midre1NQgMALRvgoykqWw4XWhGrCggvYZ6ldCuY4OOkT2/xBsoiuFL2ulh
FwxdPSg6aRxSQaLTmMaKVM6sXM2XixwG9t1niok+MrSrVxxomG47IXvBL6foU7jtV+WgPlFHmqJv
hoxMwvDvn421eFADKrMbdJCSuwO4NGHHySikZi5f+3qfQVTXB2NulCvsHgFUi58i+OZl0TiE0etg
euxyLXgqrlDQ5e15e19R0S7MbgSMwqab9Q31ZPOV7NBIEo5j58fVAQZdu1t5g4tydNUXP7e1yRiv
Z6VQ/i5eB/4Ab4PKGzdPjukGz6LBsY12rlQTbOCgCdU04lFiczWtxB+Q4WO3N1e3tlye7gH3oc+3
/jDEFclOg3IPmrTmKaktdhwKMZsbUTHslstGZCDXLfX+eaz2nTLzSQFCD4mVijosRBQ1eYSt7WKC
OLK6z9NhPiPyTkvkuilCKkLfaQC7z2S9xBy0XjzmUDmGWC6kuTPozM92mmh6ZuxQUstkfSmgT0mx
dYDaTVU/GuEy8UDELjme47DNFCVW88PPu4Z7LkDeJ7dej1tOen81zcXh7Ei7JcjGds+Z3syp+ebE
9TI4Dpx2eCJciqmHqe4VGmPoKfq+V/6xaH5Ow/IOAj6jLXuItyBSITkcVbo6U1KPxqvjvkt95r1X
S8fKTp7YUaJrqJLSNyJoExzkw7TSBycAeggLR9FNROSwpwPP2s93Sn7b/56+OOQ8lLGgBtiClY9X
xcsPGAWZHjS7HHAkSm3UtfinuMwKDG+sG2/zuCbq2qQXMVbq52ETDNaq3DqbiHlvo7VNv5u5SEnD
DGv9ODIu7jARJ8HtMtB/Ccx9W9jZj3RIfNY/ggagom9Fg7cGA6AS4z4jNpnZS+KSFAAKKzVTEJpK
dt0hzgz/dck0yFscKVypzbdFlBc2APJmnY+1RY5wVp3+bGtjpALp9mzGz6L2O1eU9OKYP/4FyPFZ
l4eSLk1rygba4nlvmgBY7I8tuVGGSh0epVS9eaLnZf9ZCZrwjDVtlAPoY13qb5HzKYm1Bavn84i9
FiM0BTzkrolZdznFW0SvRWb2xP9eBltZkD4+8JB4MwNxN81sD4/tPgnuqLB0HJ32y6Fh8BSaR8WG
owTPnNYkwsCFGlMET7Y+KOUa26PFdCgjsWbOV1DUFAziwrkpfNbF//qRrfL225hiqPuy/fjnOOml
K8ae3rV6noTsC3nXeFv/QtE3jzS7jJRgwIILVenIVZzu9tpBI4r/+0ty13rBVBlCaRLN6E/MI54E
vBk0fzsxBoFVgsqEPXcX53I/IHmK2tMUemy90ZZhS1LAnc2VH6ItfiR7ItE9IKW83K0J7D+hSwzf
WK2NFfZXbbaD9D1TkmZmdIBMbMPvsRN4IHvGV/6m7CU2ks/+clvelLkoRfQQIsvDLtl35ptAGQBO
hcBKmCXZWXCODPxEEW9E1vmIAwfmNI8ytxl/7mnWRf3ukUO9e1CUKeRbx5bRVfg43dDl5tFcalLg
CMXhQeYxld0smA2qVwmVVbSUpEJE5eM53onp9A7+VQzvBGyRAEAWDrUlQV3lyMPw8cijA4GGJdhN
XHotgCD903XyZJUtMe++fB8z7DGL/ST6ijJPTwvN+3fsJBO1ezgh43h5K6TEAx2ZZwIpzEb/+CX1
9CFxw9GobP/dpbBXOyg2qAiz3ge7pk+bOVzQDKzmTRhGjoU2Yb1W2j0j7s7gzQBRP9rKuVGiV/OL
DnQBviqH1cXDEs7Y3Ad/L9CUQFqkIybrreWZzJ+K1iFZLw33PEKKw2rla49c21Ktnc/qyn9oFGIC
pOjpj5qpkzod+qfj5tONAuP2n5Hu15mOMlMCGFjj5mrOBXiC9C6dYXNCgIn8hBv73meT1w+Np6uA
ybH7BXEgyad8x4WSDxrton4C1iAs1Bz0Hk6g6cNZW5YfodmwH48wD0sMpZtUB+yWJb91bYaF12TA
MJ8G3c9rvodgvOmb95V7v1oIbIIG5aoBqE4b9N3Qn/meSr1tPcjCH8EKGOM4el4SUhmSDjSeI10T
guVgDwAuV3gPGIIe7YV11DSYYBKGh/8VOHz4uxmm1dVRdyxDqAYfOn5zawbdoSHGUagGTOp4eEn9
hEVhyma79aqCmh9hJxmEsnPcUS+W8S3tGJfSe/h9i6v110KuReHnTyaKmiRo/LpqpfPwjpxOxgC7
zNQuDWe8y+nHdDTJseYrnxi6MxqV04ZTQy0gh6XB2hpH8doAYT4D92jp+EmF5vPKS0l5+H50KMcG
t8PlZYX6zZgs4TAk4JpLm2HQU4aybVTMhVZs5BeTxVbmgB+UcKtxHgmdp7xpIImeMkKOCIF5ITcl
5GU4hqsoE+yyCgolq+6vFwb4kb0NPr9JSWtKYBdeuvGByjPNpzbP6LQjZr5MsLqN028qn5/cKRGK
/MHPyAmz3VDoaYyrwMqS56i3fv7/UgRHn0/q4j6fT2K9J6bbPYoV2ssmQw5JWhyx5jRcpOJg+P13
FldrX/3ls0dUe6gyEydpryUCIKgx7dku+rppUa5vGIPp8cK5vuIJJIqOkD/mj+2q4VKp2DOA3R+w
dmtcEQbxYVLPWV6ashV2+S70r7PHdyQM7S4ppcw+4H1dGjOSVlt3BF3Kj4jBvdXZdE58rQwSGMlz
Vp4yTGMI3TERDLXMn8Fkl8SUQBS62so+KDGc6XvO4fk53Lodq4ScdZc4ltZcQadWxGtBBH70NcDl
zGn3Ohl7Y707qHiXMx3Cd3hkxdnBfwu9bWkVRdCFibKuEAZ+q1dSp6V4iUcTkx7qN5rIJsq/cC37
gwRelz6h7fgrWkAorD5ajZTupPIKt2TdGbejWFNpE7Iya1yX6VgEU569d8CkmlG9Yk+E9I0nAzZC
MLAKf1ziCAcckXuyaMw51erVTHiZV3hA2WXOIRfCdEYz8VGq/2jD+psWktzq8Dt6jBKoIZ+RAo8B
Kn6E1mZZeN8KDDe9jGo5QH+XCJ3FPz6wGv4Xp5qAY5bL6JkrvSLpA9+gFNHUoeU2pXBhqSQIKNyR
fiS6JhYiWRJ2e41siGFfs/Ah6OLLp/kC5rSp496OFTxRLrTXT/goT1djfj4k1qob2OsAKAjjWGsQ
ou92o1YUFD9rNwiaDhDQHQUprvAnZSTbaObeKFBwQyDMAouQT7rT8vseEsvjC7k9Rxyw6iYakmHC
lgZMSkcvIXO6YW3iuW3u+CW0Zp4Xi30ebzTPNjD8jWM33Gk4hQjS0OT/NvDFpDO1samj/mbC8uv9
ilaXD2PAHiIXrtED384bZIx3qfm4qOTdd2CNKasIhFYFxUv2nMLRwV3+wqm1MSQSS5FgRf+pl3h2
tmXJhGFM4WaM6sCYr9S0WP7jZjOiANnbIWXHky5kTxB+HObX2TixF/RupsUAdbT4aY6CMyd/coh3
ZTUYbpJSna7i5jddEmInYBzP6DU1tKi9e73zPCTu/7VrN+TJqGXNDeIm7oXPW1bh98ZPLtU2g6M5
+wvVBJlCPdcgg4s6yvWAb5ZN/Xi8jgsIpZKAvmRw5iMdRVXxlyWKPsJ8N3idyZ7AW9gb/qBnwdJ3
LwINB4Eemm6xEblrDWuCiHLp6av0qX9msduqrOgYXVq/+PYx6TXSIo1gt00VQMQ4bh0hZVXIcUeI
jK4iXLPSCuPq1bRol6EKF8XJUuTPuszqgTTlJfAGEVhSxUYpuL1ewNe32csAtM0cTjgfhSQmMOmy
AQK+Hak8iDT0uoQcuWDFduo2i1w4Z/9cr3ftXUgPu2eWwCm0U6gdJ3CH+ZX3rYvH7ly9LfXIZW/e
/GlD1AdVmI7XvOYYAZXm2j6PNfXnHsaHU8tKiKEVGRstmp+vajesLiXJCsclvJ2lDQfe6D43kYFF
cvKtGCfIH8nPDPgA7hbPAC5xaXOxqC2qWBf96UlFFXHQfcuxkM/L64Vh3D5t984bTha3GTl6Igld
X5vHWv5VP9fQWuthW3ZxIExy5u2rRF+iizFfgZYBjvh/SEYuGrZvIR2sX9/idnNz3a0k8u7/lBjQ
ESKPOHWnP09yGXGTM4MI+TStqy7GuQ2umdSCY8j9LVPXVRap+3aq32arVlG7/EWOvyjajbhWvmnV
ZofVyp+2LyfFw30pkP5M4ybG8ptCFt7SYcCII1FJbzCv2hftktckUJ7F5M2DasFtqQbQapcYk//7
xHFDvbaeAy2bUgp7lkBRNUEQkYS21pvrKGDI13If2i0WwUNzibDpnmryLKE8Qj3lQwJ4vJx2AtWt
rXXAbMg/L2NzxOjYUpdslMX5yFwTlQ3dHFAVfU/iAKvIKw24sP7KiP0e/XHFEG0YuBPGto5OuYpg
t6e24tuKjEMBzIMPUuAFWQ1FHE+e1QTaCxsXYsZovW/xry6mLTpq1WpQtYZV38eDCmN/K2KukD1k
Rz+FAxcd8ex7qjRikFH/mgl0eXnnrStfpjFWKz1dEyStxBhSpzTpB+xN9K5Rs56l3YeB4Z4KbUE+
OesGw2iHbXzd5T8RaiauF1p4RSf1WYTTa+9s7gNX66pWt9cUgfrwvRQ8z8+Y4pBz5BmPE4ZIVEXU
Ury42TasfJvKKBJkwOemSIPw+stCLZ14Pelu7shRTFmyOdJLZUpZlgZbPmzwO6dbtBxvNdQYtvW5
b8EZ5vI9oeomHRe5H7h6LeePxkckT6lZpKDgOJ7LuFJnT7AqsgUKkAwwYX8fcoVV1y6hRrqPWmJQ
CKfs0g+MvVC8Ve7+oMOjdi/ptlxWLeqmpHl6N4ZUlMOSW5arjEhS0pnolh9mz8q3ZbCCuq2rAY3U
wy+Th4wX2dkFAs+M6biWECKKLXME3Mz0jyLFwi6UQl2CTXfu8+oNpcaqcGh8x2OgTtwYtaJhj+h8
oK3EB+tvOvQXn4woRwQ3JhGprj/Pi/0Idv9DRFprA0pRK34Dxth4z0D7VRgcplY6HXvtGznPeenS
v4YVYsV5GX2eh9D24L3+/JtycMKeKuy3MMFmQO+GbiauQFq42UcsSZYPk8COPOL4WpJ4WxA7phMt
Mx1GRVn1Ac8iMeueJzVv2872BPwWg+ye6ffz1BHNfRiNKGGqotyCBKHkdMIg+rMqRZqQzENBcGRE
AHcfgwZISa2UJKVmx82Zj15RMeTxNDpxBXNFT6bjqGwKrSiz5X4uYKLVILDzdYCzD/rq0tZmNaMv
UpQHos8rCXgb0KVAJtqrRk5CxrvGEj2PsSlgGfp0RBTl3/pnZ4o6puUqeOEOF8LLfEnr5YaRSLVD
bmrMd46dRFyAY9Y7X2gI6Se7MnF+ABIoIbpuAZ1axbuXIeqLaHrOoUDKHH+XarxpNWF0rZqH2yaF
iKK3quQca5BhuxR/k/aU18bLJLK1utPh2EbBL3IdZz6rStwaoGIAkmkQctEanp282EOs44GS1xFi
RwilECD0MCACerTDBTVNEPN0t6Bf/vWcqsrdlemCjFkdKfBqam45bFHjutOtk/52+a1B/r0raa4+
g4sbGRU9NbArUL665YqMpvjJpstih9/Emq0cAx4TlAIgsa/mpD4iwgxgOfJ8U6bmOO2vsdccTUyo
+p811yJmwIUXX/dCsnKTJl1NwacbmDGott6KMvpfAHmpn4Q9PX3oI0RiEoez90I6syuBSw7xnSm2
zTwuB4A77+f7ITXtS8iQSJo2uYwvhdXx6CwG3Cm3jjPr/odVmkTbd3fk2vxy1h7Crwx9RqITdR3h
auU8LTsfuMgtd0s6RZP1YNpcnHqrjap94BQQluPaCH3TCjy8h+psvYFVHXcI9ZdPdj2t1XHCvb8A
cwy1Lnt0XYAheQFrTgCPFgpzGoy8QvKIGwERR4GKO62SLs401UdyvMtkX6+BrkE3AR8jc9NHRg+L
QXkP0iSdAf5A0Nb5NzmCF6oxGy+/gam2AqJeGRMSJe0grMG2skWBnbmA70Jf/VD5qqhJpG2ebzeX
+fabghb9pHbExCFE3QJKZHXIkozty/wQWyqy9puyTvTJx5IZdf7CCILamMBO4kaAio9LqfmR5yK2
mdUPOukq1MUVDwyeXnf0tSnV57NEw8psXOvVkMMYOiBPHee9vcz0f6hD9QRVyyap1mdF2HWnpipA
K80TF+60F/6uHx43IdY9UtDJD1EqUoKQNtFo4+Rh8Jsh+ODs9ewM3yLdf5EjJwdR0UUbuN2s+RqC
uckFUSAPX8nzF0XMVYkEzRXegKL2jtw6yowMdfeJrgkNWGE1VN1mL+DIjfgbBkonju1ZaiBGcJCQ
IlCchcNfzPddtg3DG0kz2hJVxIyn3DCcnic+aRoNiEmhroMtZ82M0RiX2o6pik5LVcRbFYzIsYJe
rS6N0H3+xZY02ptwH2OA7MmkRNuPkYLo6WslY1f7sTP+qe1B1d8khNOiD5dm9Uy6HFaGKD6zt6iH
FyTiClpyD6urlsdcniwxtafUawAJDWmPr2gkM/JyTlrqiZaWRSAQAdy6R8g1RnOpCdSzxs41l5Kr
6Qgs72ERO8kzh/iRwb2bcexYNUFHfXbY+KSYTgA89psDgqDMwrRYu/9KGbtYeWnFf7/LVzVGd+rE
/xg6AILxZnUxD1YoMsqMhjEgO7ydNrmbyoi560/2rjrx60arhLNvCFAggjZ3Ey0Vy79V4o5Cs7vB
yWxarYSYj9H+4tCqusjibpkpP7nE3KmNWnm7a7Jx6gBE4knwTjzkcReVgMxWx7DjOwRaKjL3g/Ur
gLdiGyZcXtUwZDYH/VgyTxidMUYo91ZPFZnEtXOGz3DZDax0PN4iJLipu8THzj7HNnxqUI0KtLmV
jr/pCUN1YRmYpPqZWqdu69g7+Uq5c/bs697AbccmzIaFulKuvzlsQSMbHJZt1XHUD9B8ieOTwXIE
UCRBPikpp8kDOZQOFXMOsBiY5oEHsJ8voHbiGsh5VPSnlfj9nA3Rgl62okOJEeVy00YM5cEdA4AB
f8WDA6ipDdTc2i/PMlG2R062j7YdiV3vMTdtuS7ZGuhW06RTMcRgaCwlzTp+3RoG8FOI9mc457CG
U3VDXsW8vJt2Rn1WdxVkAaRfVhi6ue0H+6AwAyih2KRg6HwrqTnx4VWA9vhK4bAZ6x725GLCI9mB
MpYJT+ePf+6y5FsUAHn6r3Cc34f7/gIaTKXNPwUVWLG/CCBj+NDd2V1Y+THHG11xUCB3ZhT+CC6w
Fy3tOvQI+k8sZ0Xa8o3TSKwY10yBo1ml0CQa8QVnilO9uaTHXg/AeMAfdqN+IHUb9oME8Sd4gyFM
Bgl4y+vXxKgfYNReRqRCmUZIrOxMvdX6C6dtNe7B03l1beVutgH5knKrUQyXxv+bB36Tz0V/nPSj
Z23vAiihfDJKXUVXjLFjV24TCkhlN8vOs1fMCRDjy+YBrss/oF1ufKpJd6t+JyBnVgtmbmLVqXlL
R7NPYLP2wF/nZHs8mOvmgsn2fFUPhAKRW2hXKI/+M5wdyAgtN5xUfOitm6UNUBr4Ohdy33y6G5zE
C3qwQ2xMElQP0HSrqN/hwglGHDB5bfY6/GWnXehUdjMn6Jnz0JbRzw+AKvNyDid/2/KfkQEgBwMj
Z1jthsIadViuil9TzjKpgf4VagSK8RjSe1ftcMXxMIPExhQIdWEtIuczn2fxPZ3YOe3EbfvLfOpv
FjjL43qAvXmCxqNjgSQUEvWHwCylj6UJthK4waacg0DfymX8Qaw0XwfTKJF3w58Htueqk8mKNXXj
cKL9UjYFnUlyWSun2fVRfNa2G/vkowVEzD3awcS657WzDPX/tXJd0G8vZpdxyo/n0KmUZHx/rAlz
i9NJlBJVONRQGYULbHP29TQxQkrVsH6a8AA+T/l4id8O/5NnDj+w/1n8jTMkpPRa0sJ1+j7siQCL
KD0siPCo/czHMHenI2gg/KxjP51TmPm0Qj43PQdgJgs485wRkrMdkKRfK2f9U93nRvo/4ZAzLK3P
PdnyXC6k+UzjZpX1AI0o2TwmwSr7BPAJqxknQQCemyFGZ7uHtxfNYh8BMXVPTsk1ZTFOklV83/YZ
k80cy3zqRMRHW+wWaM4waf0E39Uq1bb5YFNG0lJd3CC7wNPQFkjDBqwWl3cBEFrdeo+6B2HLXJTV
6A5oV1G1t9/gn+bnLNYydJ8zbtVQ4lIhEf5zGXB410rCJapQ5IOTYDCQHGIZ89dPrIFTuRzCzJD8
rIb2r33cGx6dJP1GQRXQ4IO72wHHYyyIPA8fnygffWf1+XMnVA6EGRc6C6FzhuEMqXH/YTKQJElE
0zVj1utpvJOl8zha4qzJxAgqrYY8cM9+bi3lQyqPJ2NwYY4QWZ/IpptYdba5LyaOm1n4Fyh8lUvN
cxCo2FRZPbMTyhnxjNsOm3s2uFaPbG8xYzxtPaZBU6Isn/WNG5bjlNA7kry0Be4zZZFiAo1eLzJM
r2wgEDB4RUAqCB4G1NRxdXECcaF7RvqA4MnUmp7qKH/54VF8H447AKxJirEOmF5hMSyDysNQn10F
NBBGG5lgOMy0Zi0vwzu36372Gf5AHP3l0Dxdu84uLdFegsgMTPtYtqHdnLVbHLYu2kHKK3qcdMfy
g4fAB1nmTFhamkdSVQZLjiB+LotPbz9fCcpWX7H4AX4GhiOqIgIUflyyu+B4nLHXQ60JZ+2E4WPG
WFO4XS4NegrVmxdaTDrnsixmZy+aBwsEp4479yJkA8U4FbxQ0TJ9QsUXuW+JKcypf3DJAqmRiHGR
KGJPTswX0z4QJSlcK0Odzxo9y97vCzbjlza2+LlZMTUh9xuteJMllvSWsyWPcbdXZnhXRqXGiwNF
5+x/zpLyFIVO9MrgAbl4P8wGu90jgAwIngu+9LKYxCTHwvi/xCtWTbkV5PEp/VZt8/+ebU87988u
5sG3BfC8b/OC7baaLQYloL3Gd2auDrdSJjfOSlngFEgZYUIaB7r/PkwWq4+duXm/wmxqALZmpQ/a
ZnnqwkoHOQwaBtW/mBo8ub838zMym0C8jCJ8vOWy1JZzepqlNN0ZpD6PVSyfdbcnMfkVV1uGn2Oy
g7SQeC7UVBJnfi3AM07/oRw77Ohm9evueMhgao5jZ/r7DNk3vVXEhgqP/+IUVUlyxgfZxWwt4zM/
1ieA4/roz9QZLjuMQ0HMKb90s7lp5HjL7I4CxF5P7G09vsPT4SO/oSUd+eHZl4SCZeBItVzOKmaH
IlK/BQDU1NL4f38j8QBCrh0uoBK1kH0yXJfa535N8G1YDJIjC4kDx0h47ngce2j3YvbLBe37DHW/
wkRp9ihkqC5tTs+KNQp0fNJlKqMAwNS2V12yUEcJKhqUiGQCF3iZhzSszLmkLnLvkIJqqgwqsqnK
IwopCtSIYv70n7ZbCtxZ2yh2clZ3FRQneHfCNwETBMkoUGPWr94D42lfkBuQAB5esfgLk8l4Zq5m
ZbVsxMTO7KdqMowhGZilIYrtsK50E5K7Pm2oxqwUGlivnjB46v8ql4PIVH5EIFH4gPHkfuPKfz9r
bQRDdmax+3nEwhvH9zU7YuI4YaPsbp1PbrfmilYSHyuiEs6JTiVPa7OHWJHhktkYp7l03hHo+MuO
E2Fxv/XvOzKlllm0SOE09MX0Jag567Vvx0IxE83mxyYR8IF5g112yQTArU9dTa08pWw7oG0W2DNz
52Al6/p0Vh+1tg5EqJcs2LFRhWH+hjzLRffyAYwpcFngfG2CWZm3Y62DkCRp3kUP23HC2VWX05Ra
jsb/IbKxo8ukbjxXAqk0qDp4en51HY3uYvADoog+CbLd7lwWu6aEn1N4YuX86TIHBeS872L0+lba
kpKSRiU4uj1GhL7v+7P7CaEsPx9XvWWjuVmwo8dn/AHUEmdQeq+w0XdrJJvDGG2TYImub5x1f2qg
Py92SiQNnDWYjWbIxs9DpbIxMMqS+aRBwuB1ARmV2IDRxjkX8sYlZgojrwcboaSMJZBXP14H05IH
5fUce/XpEe67vVg0ykFIzgDkYnXYsJ5KygBpPniGfKLWTZBnBSEDHlqhoeam7fWy97gpUtLoEtc5
e2Ii9zJvN+mJ3Y6bAEUaH2j5vihFFkmSA8V2fUkb4s+NpxVbbHmgLFo4FBQJhtioPlVlVZAjGLpM
KzELWrvWcIxCfrNi1E1ct5SwVE7Km6pmA/KWzqYq+UnK00LVgmALEWzimHhO+1NzGpE2ZH6TeI4C
PCVvxU9hLB2Ek/KZY6T/lf6fujE6TA7ZD0l/DKRbknWWcQ5l0VpHZEkdpZLdqq/8ttoCQh0etPce
wnFnSRaIdx34GwhLBID28zi/nF3H+pfzNmdZl+ip0q3yTRr8Bnn1A/TK1cERDagAjPYdHHXeyQbq
rO35CAmxzuB6e2etw68obVS7xdI8e/zFfyxKvo8yoZ1KpIv87r3F1lQbOVWm7B/9fnD32UGPSFfG
sV0v54FfCBG/lp2IWzVdVKzz64a7H7WDA9ol8s6M3Nk2+1YyiRFqVGEFfHgi3W5TvapvZNRSBCcu
oq6SQ0/sFCFbeZTZplZdrLZemVHxvTGCMO+DnIU2jUTtBL3aZ8sq5SiJST4Cdteu9eDpBq1SYSdv
sXKQ897VhqQbN75cC/wbHDDwSO1UoxypiM5/5OMQNRkq+uq0MuAsAnAFDSO69mCNlE1+igljZOEP
p4wiF8cX4Jz7VYThs2TFdfHI5Ig11WTxD3n/oSPd1etVN0+tNZhz7TbBE55Pdf669gWqPc2nNDUE
z3XbS9+e/5417hsw13U/p0hE38Q4U1hKEfXouU+U0kuzyZP176l+87DRwj+m0haZXDfnJvgRnD51
foeppz/Vy4/QjhrEQUmhFs47Tbo6AQt0nFx7rZ7VMHjICf+/wTXwud89mTEBYoR+ojbXPEZumpvJ
4JIJWWSiLioFIQm7I0pRpNgWxwxPTwJ0kyso+XRpDjSlJCUj+vid7TFECpG0V3IYQLn7ZrjrWmRi
ASIDxC7zgiS6EkWaJdwCjf1GFyfh1DuAz+8f41tmeXWh9klT5vGhblFH8J578DPP4CrV2ovY1V7O
6ZDYQYUAtbj3YxA3frphQsG5ld5WOvUlnMP9Fh/SRF9TMhsb5aWnrIMZ4w7rkwYJmCWhDYmkEK8V
w7/+CBw0MSdDQv0eUC05UF6gTzhBwK7npqJBd7Sep8G1h9/BQkR9zp20ilM/ZF/3pgxbRRc6GJl1
6+Y/d4kyqjeU2P3wl0ACv1JMOGFHrK8wXATikvKxTVp/Sc4+53sr77TL5i0MJR05hjo4CCOfzv+Q
QoDWHcli2gH6PBgw1bzFmnZ+GfEJVLjiHwAFGkQHuri0Q1YGKxecTrsnh1Abrnvrr04vVu7L+ADk
jxjPGxE27j9t8Qq5hBzTsG2Bjff+7qu2BxOChrDMpplheJkg3bWz7rTlCn20ZPnT488qdEgvhpC9
FRO/jMOTROxfiWYtfWAT+ycCK9SbmwdyrHQwR6ezroB5w/RpR7m+6xOyc2ip5ODPBN+L/S7JZnpc
5+IBZ1GaiYaeqBc94/kcYKfLVVSaSO5+3ILJGInO3Xti5c+3Hq8M9kNGpoIX/1EXk/WP7oD09u/Q
/DEAXVtGL4ogg8GFAjIE1vrQgkq9cOENZfC4jG1Ded/wYkZfkfbn+QmNGXHPA0Y6juIjRSKvRtgr
kdiUupDWONAJUQnWhlEokNdVVXNZURFMJZUfWdlcOGN+UBNJoMPPAO4X13NQO0bevASDl6d72gxa
Z04+YDH1Hhd7ou73fqDCITGGdNlWJLliSvvMZWpzpCAQrm/VjeYvmEmMWdew1i68iWZV9U3AskBX
TlMTZJmV4DSWbkN1gAztNnj9J+0t8pGRKo5QzzgwajWBaUy/sgr1xNniYwZi/c22erzbDIQ1KuXS
qTKUAhsDd0n6vKHWJNtFOgO8kCt+JNIKRyaewDTrl8QCdrfjrRLiNXStb9GBrN5DTdLE429R5qqR
FjPEsarPuH8p3X49MnTVLfARdA3sQbU7HI4drNLC0XH8p4vbOl0w9x8FS4fMYZd6rWWd7QD7G9zm
dKOcId6gjfXxx8eUV1Y6m7Degyt1a7eAgnIhJisjFXdyWlT8KAOgSOivtWatw556zQ6j7zduKejZ
JuF4inE/weCikz3hDeY/LD2/3wZuH9A/FVy10uK8Amcx6aUZgouXY4QfyXjdTzNo0M18GKRFw8hD
wiqPfAzCOYyEC6PWMcnvH+hsmHeY+QSTRlyO6nd/TBh139mAckIzRtjOsj2KlfR3c4qZ7YfRA1Na
QrZ7L/0uuNxwsUMbwZyBaY+/2tUNVx7lC19PGYW/fahxgbQ8gj+BXDhr04hkeUIJQ8IRv7OjEauo
C6VEsYMGkd0Va2Q66wUX6Z/7Mx6O+rOTYnYbzTFCqhtDmGFbX/oWIHr90lYtobbRW4EFcEYDohs0
a7hkuKdOI+R7IXsEskyD2bsEBSLYkGt9Uri18LxvujsbD2FABW/Lql1dITPDhonCadKt8va0lFYB
hKXsxfnW6/mcG9mewWwlyv/VJI6rikHp7F8aD6+7Cs9HjPoRZAUjeNMBo/Fs+Pik7sg7azm/Asq5
S03B6ZZKa4rUvYrSYA+jMsCX/rcu8v7PPs7RurAJi1rBxXnHwIc/sJw4BNti7AGb9syg4bZjn4Ix
RIgdkunSzJSLlsCFuW76sgcq6yOo5ux/gr8jAFMwoHb5JJwZl+wLcFvm7rXU4w29OKiirFiFgD6C
sWTHp1NIUwNvrM+ksma0DK0hsgxFbGDPGmLpZRm+p77N7APp5IHuTGorm2e1jaiz2U9R1NkYZ6Ke
n/ECXrK8atgScwNGrBmHr9zsiYHXCM5zFE7AkXGTPvcsiWIr9BTBdrtaes0GVn63AqOPHh1dzpxm
eofY7vsBDSmC5J28CbcAEqojI49jBlSlnk6/a+xHtedz0np37bF6iUtN3Rn5ZHbnbBJcX/1KJQA7
nrnqyoR0FxbWULcgamZo7vY8DA+/5SgDEn2S5JS8igJtYlyZC/om2LzwPq3sz3aOavRsLE+Rbawq
utOtitogc0l4Qz4dsrWapGhpAXSdeFymB3loqvSPa7/+6RZM8loWmnFxfgyUjc4QpgnUjsMbdDVA
+ZzCTBswx1SPNp3R1mbH3AF5V7XwpAmPtwmJX9hLfwDdbek9OjHTaJ+7L+LDObzzYMpO0NEbhmHz
tgSSyFmnUFTXVNXqITOkKVI8bw4OAc5tRjbEONpid76kJEmSdR01O3h8RQ66qalVN15F5IiB3BN8
nLn+FsXSJCqzcDGqR3fKZlwsZVcP5yummpR3iEdC1IzZD/6dgiJ/J8QEuPr5UeMlRrIUfdVjYpWP
aMVSzNz50c+wW9HV6iWANmzaZ7TTHCAWdaXF70j1fI6Gyuzlb/7t9zoxPO9EAYh5mMs4Kd4fwcZO
KGJgdad51uDSebqG//FLNQy99jAdQGahCX1UPPJ0BH+WCpdEJkKzxHYuOwEO0R7RMIkVZK8CG+6R
VkkI4lTKH8uGcw86+blxDZnQMht9o5VGnkMYy9zd0nLAQ4/evayW5fGrCMTRWUIyFqi+GUwN0ULx
QiEhwmQ/pBgODiv1cSn66dv7DvR9bMCeUsxif715Zq7BnleoKIHfy2SxECSN8csMvT8tNY7aJJK8
xuXGCDgpOPdXNwZfai2w/lmB98Ig8CHqUJ5Cgxd5hYZAivSMCbLxiheg5jMGzy5dVmG78wxGmxrG
W6L6iIzCcdjrL6irxmFklZCvdAn/exDtz5xmJ2Oncx4C6p+RoF2Fi3x73sa4fNFobK9ZL1OdPWrH
BZ78FsZT4vh1Dd/QUSTyf2KfMugKhH6xudvgURwsd4Xrxd6DDB+TbkrzRMr28rIgbQtyDyEJMVZF
/9lnV1Od6i3mbTLK+wHt47wsPa5x3TIuZbDRkVKeXxGP371oXr1oI0fgbE2kSHlUQzoq39ij+ya8
KxiNUU4vgOtefYY1boWE1r35i2NXg0o76zv1TDHDDHdPBwBrTzot8uFfdRpFwdLxyoyy+NS50lmH
uFIzf+PKUys89XGKn5GM2kHWAzXH0G1EGDtzmo2gPjHemta0rgOL95vA6AsXBHMhYYAker4tcopJ
u3+H86BYonrmDdALvvUniFa+2zSsZRERPi36o8RE7fXVudfMqDXguQfGAkR6AMrg7fuR9gjJVJ9Y
6TfFNr2zCVtHUvTTdNHZR+Xs4rzOjPyQ1SFUWoFtChk0Y/4sDRxLXjhJN/2XD1CkWya7WAW9lGSg
tqsf6ntqVieT2EEhGc5OHFkxgRtgZKvO9zI04hjnkwjnMve7ePoD/h1LZHIudy2TtAGlDw1eYZns
aDD0D1xnFrCxVb2jUE6TEIiXhM4Tb9ok0KcblCHs1FNA9GnRIhr2nNICmBjtEyfjDQA3rEshunsV
0HrgVF5dMxxyvqmiznJXZkcOkGUZPHLcOStXIb2xyRLNvfy3HDdYxo7dtZqTf/jkexvs0oad4mzg
mrnxUbHRAFbviiYcyNxJN6M6xCJH0C0nh931VRAA3ltvYcLN9whCCeFpPksrx3r4yJAlMzkC4AlJ
yA4l1VjOt3f4vcMPk2xN62KJmMI7QyNP0Qjv5kyHRgCjhT477OudTfMh7TMJy9hWu7HDrnESrWkP
HsGxYf2Vmo4n4PhWAA6RaSXScYmh7/MIdTVaZw69Iq/wLyZNzzIzLjnyTggQxk5AOqJ4uF96Afp1
0BQXhZFGQct+9a5ou2J1XcpjpnHuIAGbrCjALsNWvIDysP4Bvrzpi424JmV6j1p1eKHa44pZRS9V
U62jWLE8Rq0N+m38BEasv1kZyL+bKKDrJHLOlW2IbCTxThE2OsMW1NMabpvCl/hlAh1rQrlxh6js
7DDvoJICpLMO+eJJw3+HbHNHCxtGxZb6/vjzKALMnRhqhyiTjsXy5O3FYY+XBkRVV1OD+f5v1bCo
oZbFdFFxSsD+eQE34Y4LhrTSOjm49XKGhbtckCIFuIjRnv1T5gqADuHJmMp4ISN0E0du3AWIaG8F
8teg9Q4fXlV0U8wMDAozncsJUQ7x+IzloaTXqUdrHWq6+MFkqGyifAwhvRNdWZSMz40zZPu/soxf
1n9K+AaUrmRyPCOldRvZ+R7ejJXbSaj7Ys31LoGkb6ft4uG2kXY/bhSXQKxdy6HemXFAyvbb6bv9
vdqJVFHx09vHbi/harwZAX2xzGSkZ59DqhM61ky5ssOp6xuUzVnjKGskJHXVs2FOI0Rnmwc71jin
yyhmu3pfpZPoZBX25IXjhWqKzVShtHNjeW+AtEE1n1X0X76uMyoXt/7b9XTKsqkKOZyLCuvDWNkW
7ch6Z/MykKbfp2lWS68JKs97JEJNu0WZHcirTxXUG1V17GEL1yWkhb7PePGeH71gsyaW574Ah7oB
t213pGIvJ9acyX89VMDA7uxyk5M6LyQqedKuY8+Jbi0ZlO2YthVnYZ9AmW1xo4OQXAmR+3QCbmXV
dHi7cpEBYvumOZelObKpmXx5SKUh8NAn7j6LjpOJp3sZmGFPRE5HA/+EIfTsaWaJFG+rGosPTZYN
GKSWaBvkKeroechiblisZkVY+wsQFgCm5lEn7KxWB1KfqCRgH37laTbp8qINLS4L2dnEcA+16Gc/
l6vsJMbDeO40QNyZAq64pKlAMrln0ITHMQfDValrtpUs7f9F9bgoi/IY6sVuxe2LgLwO/A6ftzTR
JW0pHtvy27lboTBHpXLk5NbHbp/JDkE7NsK3Ow7/qwGDknCmH5k6FKBHOum5SsRqJg2KWvHAiQf1
c7Gt80yUrwsRUUKpRFQG7ekZpPhK5QPEYj/0HaBiW9kU3WxCXbJCUnPxZ7dfL5+44Vg70TLhEgwZ
8bYnP9ijPnngqme8vSXLwCeINGuS2ENjD/fJwvGGJjBzXSGDSMtW275gYuQbHfWISwBcmslQbtah
5LXgaDHFK/K35eigtvC9ooCkJGye4qrE+A1vtM7bkIynsfmQvPJ6RWQNK2nQkS+YetcjU+0heVwH
RsA0AP1DVdNOyiTX3NzUME/qPPSmqQpGAbG92LH7+f34DqFzflvPtZREJ+ANofWJTcs+hj6O7dHv
WSawS+WakfZ2Q5Tlel7r8jfy1W+/nu4u8RfHn0Qt3KppMtnqRCP6uRE+X1/fIo1cI3y6vzHCm2cF
+dcEQMrIAQhJz1e+gxcG4Gsifw31zynxnGdjv3mT+K+WMbEHhGkqD4AI+eOfy7po9SJoCODeJeN6
z/Hs0qnrDpRGBEFII7KG9U1rapzySfxpBupzwXaxu9c5A9ZOqQRQYaDIuZojME/KPjIykYY7i2i5
jNsEy1frUP0l8c0kG1kHE7/H6ZAndpJ+Q2J0VTWGypOKOzmIvKyb7oIAtr+N/9dioWrNOJg/dvSi
SGsIeKF69vtV7MofYNaw8tf/0D/B6w3fh4L6aOR9qVE0kHxr4Ifue9ir3Lo+KvVM/AyJrY7Jmm/P
hRV2jsgFD9pPHULG2oMAubXFagqH+vzMhDtEo7i3t7xqEOqTMJgbFE4BoDfDOLeWoay2Tssfyipb
+v5ZKmKNYvliHxOXd9KCfvl79ln1Rqzh8nuspspY8lvuwCd+UpVne+9KS1Xj62lwAavLgZtbsyz2
E7DRUzoU+c+6pI21OrFploRd5iQsbdJ8KnsjoQpgkPhNJCa1wqxef/2+5RkkNtuN8lY0vfFWdgPR
jIqnHvaGVPWQaTmzyWHc0KddKp1tKwvJQMq2ovPWqcKuujzBbE4zTMavNC3Vd1nIO+NLBVkAdd5p
JtPELXJklp+mUaYbpAbo7PpWBaNaZeHt7/ji34aoqPvUlg5WkcFl5f0bWPwxJ6EKYH9EOprS53kM
BaECiLqXlDj1flfAmEkHokb6cVsCtA+7SDOO6fuzuZKAnUI2ehwjE0+WK3CrhZKYMn6stnQIp0/v
BYs4cTNj0k8yz938OjZxGfO0yVtRcsSdDwz3c04P5/ChioVcqHyuDfIH19QSycXPiD/IfZWFe6b8
PY7BwQiVFAzsy5biaFzQ+pqP/3WxTgxXyySgaX9AoNqwJIaEUpnRrT+iV4lfX9+QUvqK5hHiEict
58TVknhBcWB7GXx2f0At0pYDmY+6MapRRDgT58AGqKF2p+Z06Xi8fHw2acZETzOpJUkvChFBNp97
eR0SATDX4/JOOxacNhPvEhZKgVVb4ToaY+0GguYvlPjuXeldcTFMoTdhjajk4N+sPAuMqI79CVHP
IhZK/p/oJ46clNl4lXxc0YH5PaewDwRIRDoeM5U5pJEpJKOWgwOiwhRFX8uGNBXy8b81XiPq83v4
nKxeUGqNqXOnJwbsFo3ZXDYj6QTzVA9GLnuispqsltjU+ImkSxZp5blXQDQecKXOcDROCGllRtq0
5Cf38mV3mlw9He9OyJ82mhH7W57EVxEvaepOg+Q1Ufr49ORt06DPddiV9lWVE4c5pLHe9CIcHdfs
Y315U9J1VQR/sRuGcOOYBL9Nb3MEyt47ZwvO2oOhu2tGJNw9NhbtOmru0EdoP/w42CVktXPnwpQ1
CVqC1ywGjHijesjcnScajhPSLf059/tH6q13lgG7kXRzlIdAhfO7zMtn/8xRmlxjKQEtnYlxESiz
8sLoOPEq0mz2hwl2SL9WtCkvcypcfy3wZRksWY3U6+LGTzup4UZ+SMI4W23Fxcg35L88mQmLfTWV
IGKJTXCP62nzmBLMN2tN6oqDyc4BvQfXTvp4Ca27acd46Wti/cH8nyURS3I40XX11Ad/rbNpt+iJ
0oGyXOd9ViKJLICG3O6bnfw4fS450FftjhQf32Cm+67/RBDFjceOrzGywcOz+uKPwgmo8Xmq/2WB
LLVaQVkYyHo+iO7/D4Ii2v2qqmhAj6AghhJ4ULnidexe3S2dn3h4Iecu4upD6+kZYmK/mDYmIYpo
cY8dIxEmsRq/6IiaU5Cwj/fFSDxj5yNURYTzrzze1yBY8W5aKG0s/dJ1qqZccXzUl2tfNFcJuWM6
MPPq9BbQY6/YSx99VFYjXleMmy0KliW1NS8Ro4RjsZP6sloUq9ndsVGpAVHPbweyHypJiCmxKE1g
9WmRPEW9iqSsG57GIvxheCvndpw8u91n8bD7F4QVuVIeEeH45K2+cA3s6HeQWjOhWKS5GO0E0N5Z
Q13lCn/VRUEDwRMHQg/LvI9zjiO85xE76ytjgQJUsW35dGfivNOejMFEjn9NFteqFZ36mgKy+pX/
IVnH8rr0uRKcpEXMNkKCHwenSgroj8mP2I0CMyc0xJkY5V+V30HCbcrGAyT/R/3g82efxyrGqQSa
dU/RODsid1jkY/yaQE3W0LVC9tjlZHU9s/HIxCXkPl5kHCny+vny5EWDfoQdG5+u/D9Bu7DlC4kL
dVcgS6D5DVdfJ9/cCO8nLrhrmwQmE9G+j44RsboWr6M/HRo+dqk4lPAKdfWIB0uVsk1DNXaX9s0W
LFDHmSNr3PPIV6FN1uYHQuKFs0Vo+BPtVwxHs/V35CxLp9BIwGZmj5hESrDhlG4iiij5H0E1WqQR
/qQ96PFmiMcZS8OKnbz7WlxFSJEcdF8V4Y9Y8yFtqsFvux4WiGLjqrRUljx4L7LSn4DCMq+g35us
rjqSGb9ZOsOmPb5CY+dqEsz+CsDwt2S9LgLs08VZsu4mGwSnh4+Frm9HEN304SC7h1qHWr8KTJpA
o1FHqDpJZLvVukRRfgRmP37m5Zt8kjvLSx2PRgR1ptlNcpy/MdIn6/prjFMBN6UgWx+vXmGwuUPF
HUx9PXsAeyfJGor7mzVo0exjQoC0FaMuRAk3U288KEGr7CPO/CtBjbIR+51yQsOK7ppUPvuURKUy
AjIveYHJqnoA8AK49SYIRJh24ukEoWXI/T5vHF9oTzIRJvckQdeGBZ3q1l0A1stPcLtCiqpYtdA/
EpXMmu4uxXE0Y9KbnWHGGPHdsv8pIzx6oi5o3nJOOMXVOCwx3jbUk3JXkZGuX4B396E4i9OGguJU
ZCQyv3FYw9I6MGuGTFGFt0cEvO4R9w/qKh6Ar+IoxPmp/pb90qIOBky6bCCdS4kbyq5hpZISXRVi
q/aWNregh3VYegPwht68n1nqtv7Qy+mGxZbHU4QxXG8BgjHuxCGQySnEIfA++atrZH5xF2O2GeRV
j3ouMd6uRthcWKjJumUlPEBUnl2NssMI1cARRSjFXbIEae/Y/siel4kCdJG0R1ruP0LqTXqCpRGN
UUGTdCg1qQB9lpTV+pC2iB7qbvYYFqe/BLg6ZbqwgZpvczaYjM3XK7xRvt4Q+9cSoHg3Jey2qxCx
zFGWP835WweHfV6Aui2dUQUcGi3pA2M2EUd65afSoUDtsWIMZCMBqznZL9aV2ogo2mbSVOzQiAMK
mhAAmzTlq5hTpHdgMqpJzz/X1idmI2XVTpu7AKbaoR52usHYGXw8g1VpvvNnpaPjkAdIav6pla61
fHN35SlXnc39ZlUjBkcBWqJjgp1wVLSLvj4hl5EY2JmMLPcnUA0uymq2A+sjUQY73hkBQEzgiJAp
h8SDQoqicBorSnr9aXOxar5gzoWZjjb2CmaiKwhftobQqwlhW/rL7lUQoT6264vRAs9fto29hDqv
Y3aPRUINjkTySsWL1/YEvqhDJ96plJCilG+3EfI6OKMxPQYpSHUWElL5I+4A9Ne4v5DKFz6gFbAw
mPW3GKF4NWbG46eL7daxM8S3kA4L8++gGapoqRFq7JtQaoBPg5MKEzUW54a2WoVfzn2SNLBklYnl
f1cUCT9lACoO2eMve7fJHh/v8sLbTe3XzibaPtU0G0PwVR/tTBGiZ0IT+Wyqi/KftTObCJSAitr+
iMTK0FJXA1xbcTRNH471Ow9bw6/tVQA9LzyIPg7tuWGY8JkLMv3p20KNYRfEzyDk5v0PgBOaAVk5
iP9UjdBSbwo1gGulI30zRgxaASQjDftN/wwvEqRrkuV9SqWHrme1pVKHhRZdl6jZyHHWxuFErUFb
1Q7paGuE8xhdAZ9CUhP3UNv8Ope35wU/HKeXzuaSrPdkhdtqIChhoHRattcf8gOGvJlG2jNK2Vwt
uDiHadNhe+7asbbJuY6L9xvoqGt5jhuqM4ep+7k4qxYDTEwBTA+/wFFXxqPHwEka4wnQekyZqwn2
iMYXatptHC8SsY0WVn6+fIn3MabcC9uCDSs5/Q5Jbm/CDD8lLLdwDQDRL+wHlpuIuOZgnvej79zD
zVj5H5g0oPqiy+4HzDAsDaa84r5lUuzlgA7fmoevtzIPnDsVHV6UjIPp6Kdv4zNSp89oM1CzWp5L
lPZR3AI/pjVQSqAmzzciMIdYHixuRS7EmqTFVq9srjNuuaCWP3GHtPUJA5Sa1Iwl7rmgsFtgU4r3
4bAgKXi0gy0SACTK2gcPddFhxfdvbKa1qQq+zYw4ko1UApAa5phiVae8sm8eZv5+D6TBBkUlw5l2
yHD1Kr55XXcTTwNPEw9rMuGHFqxSpxocqNAmfwIDrFtXECd8EwgUQyXZoEAS1k0ezvWsgLxxJZGc
SjCgW0eKVgxffVGou52fvfqywb0dM9YOJGNXPY8eWaFYs2gE0UIZDrunqhpALxZUj0v3IiUcA5GP
FRY3GPOfQUwTDBRMkmb9m1b4o97sfmMJfL0GOOKc4uIcN7oij9k6+9wDC3ex4GBmunS9NkYXdivl
mmw3OMW620jWggisDOM0KhfTCBYBy44O87M8+GJBMjwRqI1nVEHCe0sYAnRVl3+fAEIOQTuwJocy
62RBbdDvpisJ3DN9FH2RDg2guoR1uMaZrRFkczS5LtaDVaD0MuTgWaVwIbetOBLvq0zr4c0a6kf5
HeYVD3P5tM6s9SK4ZZIsKpQ8CRbSUue1hIuGdPxe/P6QOf9EUY9RwXe5k5Q8lkuRQ++00Jqg4AFG
bXZcLxF0NdQuBxZH9FvWSSSSur4D5LEX5f6cioBD8AHeWNwoEa3f3xH53QLXIT00y1soVcxNPg9X
luH8FjO4PBkU2E7QrZ8AMYsukPISLgQXUVueXTEagtq0PNgxU9L/SF/4jvlqvMUM2J4Ap/YtJBwG
O/qHOMBZ7Z66QCveo6G5wvbptWVrOJIAEcFazhFl0LlSkh+iHIVGSgVsGLdzE8WTo7TcJrDOeMQV
c01JbEl8Oyh4jJ9wwlCp3JRJ8iDektlcZgzuCGjUAC9m42QdTDTShG5czVozqGQDjVz9sH/fZZa0
CD7JQAD9dQ0WuRuzRI0XMMdffVePJDGucf1RTvL3SLqwJ8mZU07ZC5UAwbyxHAmZ2ENlYN0Odfgb
EF0ifjdB/VYxcmcRyFEQ1kf9Hx8+/vKrs91wUyi8ei/i//J4FNgwFXZMJJOCChAGduGfgX9XLdMX
gg4r9h7oMWE1LDRkHIcseXucRS7g2gqhGON3efnOq4lp4wrPrl43zx2YsJzIHzq4FtQe2WPRQlzs
8G4XDzWiwuDGj7Rt6Co1ShL776kJxom4mLmkH733NB4EmsyR7Mp5cZENLsP+HwGKnD3//PtilPqi
1HplA1rsmDEp5U+mijpQT2PZiwdh8aDvXB87JkwWXhuUYTh1Xv4aCOF+oYu8dONSkh9EAwLnNjuB
AzO+js3KsrLU8BiuAtHFmQXTSv7hmhQNXjsKW+zpfYICT/DHPuZfp65qMSkZVoanf7Q5S8jbiRxK
dOSYD7hcNnSMtjwNUg8HHbwenoljunT9QaNfKo/X7HabwOqVXF2WEydWhnY6dHRgIVPfmlpxL+Zf
ct6tU1Mg8bt/Ijcfbk2vjlk+gnQ/+N5vEa8z2jUra+7pPyII0w6Nhdc8UP87m2iAKtraX+8fMvV2
PZuR3h7pEND7aJyRBQsz1I3937eGGr0ctt6tT8fTsGMs7o5Gou3aZxtSU5PJ9n1ExAtnVcD6Z5Iz
zrH7ffo1fGjxmKZ7/rBJDxGA50dG3KJdHsJ+SsCAzy/gfX0ASMCupuTeCsXTR/ty5D1hzEeMx/ns
BkosiuKeCmE9r5NoRuBNKD7osR5gFkXv1+5FCmsGKS+D1dcJIncYJCSwaxQHwyMrDs2SgXf0X9VF
51XKXuiP0nT8Kr4gsSnjp7FMceTjgWACJl7ZHOWWi23Spqcv7sfHeHanavwK+7IrRtTi9jaxfXOF
CImKV8Ea+409jyLZr1cI3ahO7wL0ooK/zERJWgk75N1wJKc5RV3ZGFev7Umi5Xj9fI76tigXKz2x
4FU6NWFq+DLZQHwq77aJSULt1nVesr816Cd8p6+RaqLjrc8rBBOfTEKeNIJz4KpeWMXCVNIvHs/w
wf1rtUkFp5f1E0O5vqGh/K0qF+v7cxXUdtJtvPPV75HDHdrM5xs+T2O9E+boW1D5YaFF7sHr2Q7G
MMJ7gPe98hxdkbLdWuuAhVCRvhfPFaEK7p0vDY7oBs1Qd8K03bi0qjLQkm/DSvxc6zoQ5pZRfqlx
Pz/SWvhITtb8fLF3O8IE/fNMWX0k/XY30+e+6HUFmXknbsm5KSWg5gUAcy7OIqMWrkSbXxoX+1lV
poWfBCJH4JQv82wCUNUxM4BdJBbPOdZGlN39wo9Q8E1Xv9VLaePB0bZ0yrFEDTa905eU+Mdlq+vp
7dbE844ig3rMV7zn6VchSHiBYVAPdv2vgnQaFIC/zEGKyiRkVejGRy3Wdh7G+w9M/eIGnR1deHvZ
y+DWP6M1bBRgQDTh18zBPIvMbTcbW9R/aQGJNtoSwyrteeR1EkiUjpelu+PHF3wuqlYluTxGM9Ue
y4qGYhZ1xlX01Fl/iVnigAMgXEZ4lIQX4cHO7W2UNKQ5ClTgKAa35zUclVG5fGXkwK23zscinlx+
ZkXmrTtGqPzxQF2dv7c/emakawRqq2c3xQqGza+1ATdL1DoargsUO+mxMvyTP+5FQ7eOYCotw0PF
dJCV6lKdKtxzpOtqtG23kSM1NHWyq4qgSIgyD/i3/Dxmmf13VyZvdSbs7m4YRhnqhNASps/OkCuJ
YB6mSWC9nVhazKCLQBIqZfL3VHLuTe1TCuN8q3lbsgez6LKtDjmvWKbUOcRewdBsUp3K5Fi5X4sw
fvE3cCgTFWaJDpSf+OtR55osGyDOyC+MrTE9gFNv8aXcg9xVrEvXTiUOCXMjsFpfpKDzIJV5khkK
OcwTuTh0B+MGn6QGf6fArqSVQGbT01CJk6beAe2KWMRUMXJwsTb6x/nGixsN4vRApMHg1YSdKj+D
f91F8FergSYgkbYiiGHXZGB/Vlh7/KzaXjx5MLd8LuhKY24azBlPFek71BxexAUsWiMJ8lWLVvnJ
V0Vc+mlFZJfNa+XuikmwuD0ZU+TaVkT7BkRLOtL9v2T5Z2gx0sSG4O7SGEu5dgDYl4pR8NuvZRKV
ahGtOxaBVHuT5d6WPw+Eqf/MHMDjTEnpIY8WQCmYZMsipkFXZmbmXGyrsRu97/v5GX3z1iHpTacb
a74EbZ4tg4A626Rz5ObxkEK1lMpjyqchT9knZrpgIUY6PhRlEf85hBQa0SEpisysmXpjQfdFw3c4
NVEYeARfP3B1G+JhhXwKO0MegVzxHYdPFsnXqQgIJcGttvSyPgMm91HsVbvX0DPxNQ5/DwyXICav
BnCUOQW0hwW90sTX9UXxjjZ8da7+i2c0uk4Z6GwIwLP14X/AzlR9IZQuRdV/T/SvkTdECs1wBKyl
+YTf3bUvTj6U7zBpHZaPPrhYXLQhAA+e7KRX2hZdjtphkFkdURDNZqyTUcSZiCsnkX72KJzJI7R7
omJwr/vdX/WtHqRJX2ZM7tj81Ghfv7y/Q9AfeJD2u2aKL3kfqzkBMOq8/vRmNJEdBqzoIh/SzHOB
TB3yhLg7UA1lnKrj2Z1PEgabsvE72v/C/eZ/ubYnLVtR2fYm4mDRnI5KDPDpNdvjtLu7LTZVP8tT
1f4dauYxUuPGZK5phCiol0c29YVRxOnl3Yx17L2txKUQoknKcE9tqwK8BMr7z7lRj8CCaPAuAqz2
NDpTIfJqU0AIOVfDW3SN3PE9ir2SJgLvqspDVs0sSygoyt+V9cMdJx2pyq2SybLPG6UuX1UjOEng
QiRmyvnE55Wf1ZP9Dje7B4iVhtkDB8HSh57yseY7zYk8gr/J4cYQOuWN05Yb5wLd3fFQb/Iq6dXR
rgHPS9M9ia00oiY4QsDPp+v+M3GLc9zVgMze+6fM9b0K+V273YZYf57XORDMyau7KCFYMfLMth4l
L854T8yCLK+ixK4o7LPEY1A4kK+WpgbOowv/lH89fEM2oJzbD9UFvEzf1mq3yhmDeO7hWZRINuTD
olUAx1xPIZyjIsL0zWVE5ZWbY9bFbfCSDxB31ofhQfHpjXT3uYdOisL6itUE+NqWayMr485Ec3Ei
aIwnZVS/TwGO8vUTb0/HPej/0iHJWSH0sXyR4xh0djiHZ5+DJAcYTNjEeRR3oq7NTj6gzH9lNG/g
iCIxhAI2gebbJn332fw9In5x2JV7k+TqULY4mj23sLKOX2wdV4o7LME2nrNWTIrtVHNoBiXC8vc/
HkuVM8HvlCVPoFATXszyCiZf99geVy2XGOxv3M8dJtw4X6UG/qkCsQWtWN50ROCFq++fnv8fldEJ
1H6ghbr57LXaytwd+wojNHtILsRDePlCQfiTFQA4zK5/jmqnDDm5g7VaczYdBZeWzwz3K43ZvE0p
al3N1O8DN7x7ns2Pnt4KYE4A1omDk9igxh9bs5PsJYtDo7XlPC0ZRS2NXLOh8+EwHcRT1R+EAy8O
2jekco026zl85dzbb4SS2Ta+DvF/gHaVd+dOOj3F9rRLkr6x7mwy7yDsRvZx1K1KcIljgm8SozlY
WD3NAuDg0OsUX6ysFfYV0hMc8ppF2MU2+AcjrFseTUP4XsKWEmktcqmN49ftEWYwj94+B0u4SI2E
2ssmwkQMb2rpPAirmJvRKocMptsvePdSBJFkGVq9ZfBzBut4Yf4FkHM51gsxe8ySjA1JSB8hmTNg
RNVxk3j5RLfALUKvbu44kDYCn7FSOOsARus6y3Z9xu5ns9t+s+4pHcdJdOf8fRYHjPG5uo0RFW4Q
+f9VTCnOBHrqx9iJnJyP2hOrbfAY/arJc+dkDAE2apEl3sIxZpWW8kNpiCSaE8N6w2grZgShPPuN
etJOOSnZnsYufVFcmrAEC7ex31Yv6K6+8GIXaPPgXX4L8xtQ1IQnyozmeokjHMxnk9b2vBJ4Ozs3
l4jx2f8VK7/l7dx30ylaet0I3cOHOtrdzsbmldCyMxp0KKCczTrKWcNpTjldj0JAYVzjymL0KYEt
nEKcfl9YsZzQhCIDBITkvsfBwZEqT8aYZocrLa7k/I3VHJIYDpQ7No7lZP3n9IX89V+EAi2lDiZe
iCH4V59sUahEOlYU1EtMgd2+fbWcc8APDLkJZ65w8JZyTNJhDRnM5TBwpAduvX+zP76kLSSaez3P
HRkMAEw6s7gL0oRwPqy3MKCnNT+C2x7hv8eHQcQoa+1qaOw+6Z109+TWHGrZCkxSUsmbGZuQsgDV
bpeYpRtCc1pb9TOOvUnOPaGElLyWGvV3SIRS9PDsTTRWBcRE6RnEVdMeBRIUvYd2n4iOxRcURgdi
de574dx4NWKw3je7KPZQjvBu+pX9Yn7DbZr51ltfqAMZcdUd6TwFtiT8njUq6VNZy60ymVyilpTq
kTbKsTn/I+gIlgot3eYL9MwZV5nB0rgb+epcGJ+VTdF+3hcxo1wOdyz927fEkPBQVkqxLrFZj2Vw
GGGD//rhqfrhj7stAxwu4Cr2JvaHnBXoLZ3WW7Q6RB8VVisImAKnjMaA0S0BH3kmj9nMxM4Ujr4R
1Pje5t8dmc8/9OJCeyJM95BKOMfBpGANTeRjjKJFTiROF1RxFNVBoezvnzj/Wdq/IA5MhH9XmvYR
jqiq3MqpZcJ+/yqi1zQZbVXTawOcwv/xReZ3bG+sH4fTiPsosVo9Kjbe7Sr5Lip7A+dwAPtHEN6u
QqK3oKmrwdv7QddjrsgPXINuH+1uykcpGwgQKTyd+PWPXtJC3onOa4S6X/KqKpUa0Aou3HsRFodI
TbrSMIRlxutB8jPCOLGbuMN9JwuDUX8qv6sw+WNbSuhXDU844+k907Ts1meYgn894C7jyM1dG7xQ
DHArty9WABdLDw3OGycfyLiT4vj91UIrcTo1Bf9mQgXkZUkghgDXKqztCWeGSSz4VYVeXtiY6qFB
9QS0Y0nCrbcbzatXir2V9PpsjsL46nLFbXj5k6nWdYioPc2oz1GTmwb8EA8Ax7tkFJoPovoyxndK
nnQQWFZOaNWxnkPLsPGU9Q2w4vGK83lfOhxLvAXrc2CHFDmdlak0Z4zSzJ1M9V0HMygfIRa2d9ZI
PHWVK67vdIoUmiAvoiN00pigbIqiQupUgQi83eJ0OWUi1qyM2UhwyoZMvmdCN+4WqhzmbAS8tQrN
vIZ6cn3NbFY3kyFk5c3wrPxikvpFY9xKPj4EfA0XZXTr2s/CEpUgsUH4afkUciQp6/GVzZj9XD3Q
A0YGymztcygfEWbNlyaYbpoft5gw1RAHdcVLvkc220F9z0Hw2v1cgeDTFkWTUw9+/4z/l/prIcjA
9BsljcbqBF2/qxz7ELHzxHXctgIQKF8cim740ZxGOYgRH21AcOfA7TTuI55YQiIWx7n6n/MqU/vh
9De07gnsvWJpKfv9JMSwb/IRKC8Aklk6o/KUkG+E1VvnCgve5ysQzFWNtqa7uvdeLivEfjIZtDvS
RPdJseksGwxB4IJoSP7m7Y3/DdVP8o5WXMct9ZSzngKu0yw/ZDVcrnXFiRviiigVSZ1TDErI6/Iv
YAVu78uv5uVjdQBU6cAD/YiAYn124wdkjD215Q+ofDOh+2iD8vmRYjUA9d2TjMEF7i5EuXi/Mv7D
0CwXc1neaO/NlMvz4pVWvu6Y5fJiZ6v2NW9MhGkDB7W23tLlSIBcQ+wd27//rhSZobiIyRyT5R8g
W79ZWD8jc5tyjMAPCU4HESFIlZ1w1XuGI+A/XVqwJ+nz71iHm8dteK0jjmQ7eKp/QavdgrPgiHLu
cpGNfNIP7pdjLKQrFfy6PUhEBL0it8KGRZq9xcqKsssmhBP7YlMNicVPRZGjlKb6g431+/ThGppq
UbUQgm+JGHl8L7UqQPV6P9metN+ESxS9mUF1GRsLssVCfu2Lub87+HTxlFnJAW62EIFUhT2rRq26
KJWnFzp7nLzkQsbUgCSjNcB9qseazjhIDz6MkZoI6xoUVfL3sG9pBmvzp+kelYAJ3SDwcT+CDEzI
FCZHrvzT+Rw+VwlQT2Zc23cZJAyOj7R6jj/CeyDaXnvAqdC2aiFFBBk8I+Ao593/4NhuRivlqK25
1xB6cPvroqMMiw5BztUY8Eh9SLqoHyeuVnqfCLEBtNCbtLsY1euNRag3qGevLofK30gf/URKymzD
zy4k4KhtaFkoNb1g5erfjejgQNyn2SiGNltQUGOll1ZNAqD6F0vOh5mAclLTqmJf3f+Iv2T0xtKG
Ml77LUCVxajLp9aIPUmYqG9B1Ttom7aFY3AerGWL0BPZnD4LTyuCEWR1RYZAxGR47bWDT8wDWyQg
JnFmpECMUZptjeTZ2S351rAzJhZR0wNYH9Er7U/YlIcoacVe9cF9qV4s1DXtmyzPm5WDpn15KgbT
YZmphlx+0neCu5XMTMRu6s0QSmJ+zMiQ5+JtLt0470dla4pXblyOM+tcwiSWic4775VSUTZWJYZI
Ig5edsOtDxWn8J5Sm8iRUu3ioUC3AQbz6PI9T9mGGrxuLw5dpwNielR6Jj1Fcn9/MsCJSMdH4DR/
emvDrbpb6sRmOBcU6y2+6/JEovUgYnS15FBlg8RZ61c6N7BiRdRm+LSu0Yx5Ip2WyOyR6ZjLdu/W
Y3p46LC1rGuAkah+TW55AfSM7zjXmXvoDVNCEgNRBaMooSKlOGMUwVtNl+q0HlGWVVgcqyBVEw0Q
MJtlB8MujSwoOVPJq7mjTb23cGEu7x9tstw1C0ajT5Ic8yCAaYfLO/c+xxIq1NeVDG9hCEvqKgXY
FkkPNzVxcxFPJQI1DSbCEEBjsrdygILgHy1jLnDw2sI0bb7nr0GoaZWsA3g9LyBdrvmbHixPWUvo
IfDGjlPV8UGNdTYa+oAh3TBWhV7kgDUvQhgoqVbn1nUgmCpAo3xVdjJsa0SBdDuRBpCY7Cm9lOqK
G02ZyM5kQF5QCgy6Mzr3IGbfGbu+S3mbSNBs+L3AJYgcoYPfa8JGG1B3BJ9cZIkALbbVzGc9GWjb
j9LI+dsDFgkZa9hnjTO5GB4nYYTAmmjLoT31exOJePIv/xqaHNMXItDzB9gWO3zvJJB268zUlofH
Mc9HEN5gYzK3LK39aVszKinoceH47RCQCVvbsqDl/XSIGSFC4MhwullQhwFY+uF8/dOEVOy/bkNm
skIFBwwa7kvjYo/HEx5ALBbGBkTKzq6Xsxm22ahVw0IH2hmiBt8GmfDzpMcWJ/ixBCnEym01czAp
mKp27L0VwmEjv6vRRNRy78BmAUWyLEVRaEEbUs5Ty1gnjHzavcE9mFzGMe1OQzj0qLCRt/A8JosZ
E9lygTovjtwpjEpZu6OPKcu895w8e2w28TkxAFuhCW3njl+DJUCV0y5geCiJMnxYCVw6v5s0Dfx8
w9gVRXcKOXV9rRX/7CgPcUdjoK0EcuFpFep82b6KKNQpE66vmyL0FdU6gkS3z2ASMfPpvKkKwdhW
fF8Y1hkJDcyu/w9HAAv+dirl9gMhz+lSeyTQfDYitfaYJGhKdmw3U3Q2zqg8lDKDNIOhPCUkCeM8
pOIrfpuQAR2ehlB8/clCXkbnNVLVBgVXNk89rh+KXxGiT2adOc0fN7oJkAKN+/DW4BJjSkDcuPOe
n6POA/K4eNHOWjZxuGuFsUy940svlFcdmLLpBMdVJDgtkaEAcXM5aPb+gnaxIB8w/KsAwyzqV6Gg
Hhx1f6N/Gu8b5ZKbOfxCbBlr/WgFp0lZAoK1T8rViilcprydAVJVXGWejg9mndX275zffZKh0Iwd
ewGoMZgvjoowT362YUJHoMP8PEfJnQRd+R/RIUWTsYYvynq+QppyqIJPjjldawmP2AqKmLTH79DQ
yV5APSt+OCwCP/pEu0RJ1n4hAqlK0SW9kmPAWbEgmzq27tUcIsaEosjuN7iBGCP3EEkhO5ubUWDK
YpwFiz8UYjsFclbooXCyXw+fg0+IDFaVVdx1NIv2+nxvSdBBFSHOrKZp1EzX9jzG3tvGiK0WjHuF
8VUFXh9XxVSM2oavdFu3mN2AGDfrnyl58wUKJquPWxHW1J5EH06XPS/6obODMLsG7ZXWm6Gehygl
X6No/vn76oB5fln18n0WL2bOKKQIUisdRizTT3T42L8fXPlXwJiu8+JOFMGZVnjCEbpUjaTHxIgc
wxrEF7zAVCEYnkAg1xYpAAdpNwBp7DpZU2viE6iLsfgjCkNaEHb1Vgd6x46jCslHZiq7Yxhve9QT
4SFqF3/sAm0VHWwg8hjKynaKueoI/R74yyDGK2I4KhrI4zDWLpwDZzIGGti8LN/EoBdmb3k+E2yB
R5hzUVP98hpVXT4VRgdaX7gqOt5KX20b+2k+ZDkbdv2DPLZMlWbI0qJM5Ygsmj9v2UMggQKEtjNU
w7pSwemvI4aL2M1qmHY3a5OrxNiZeyQXcSjfYPyUfSNCInyfJll9HIXY5fYD9k/lq8gDojoMOrKD
J0WutdOM85UkGdMaTB4B/msJQHg7Tcmr5YS9XCi8FavQkggy8ybquavKFY1QoZm+N+qJIrS2K6OF
lcmjhx00U/mJmwLCykWdQsK03++wVkv/31tp0Xa9EgMqycNZqk6W3dbojQrKRgmJQKmYUCleilxu
TS+ua50RuX0F5KJyinLb0/QmMdeLogydhQQEz6WE0jlVQ9DH+9sKq2H5Tn/YiLy/lMayaqSehxbd
zjH9i5ZdGI0PIp4+wBtKrXsvAYjGDzEOFwgF+MQ/ImjTvQtMKt2xb+JoZC66bnsGfI842qDnj6AM
seUurQiPZudh19kPxqM3CNaOi4BWHs6vANm1x479lfNNc9QJN1AsJadBeY8mftSAsY4y3FkMSSbm
nwRBomiElJyaT0sHUjsJjk0ILTSnWR3QYA+n3vdU88PLJpF0iBloRrwxaTS01hphcLEuzXoW2AHT
zHPFUK+I9BtghedYVG6JK9k8bCHGs4CsGmANedm09x4y35RqDOQ85lj5iQfEeiOsBLmaZtQJStps
2k2HSTHYfDGHX1+JsF1l3V9bdcuvIGiSBsgCq0/C1cy12Wesqfa/eVsH2OdwXpF4NjEUwsgTdxA4
cumYI0vXz08eMNah6YqmYYej51tkTVBhEcPb3GIQJoBwDrL0UFPWi5NTLKXceD6DZxT0VKQzPT75
FcPjC8Z1IR7m3FG14iqLF7VlmXszMTfmzDwoJ7wcT2vJ3ffMoCyo7cG/MUjc18Le/e+FuVPwFvr1
3FJVfFpyL4aWMXF9s3Nl1AwNBa1NaSjX6prweu5uuwDiT+qK/mSNX/bkAQZGHjItJ901oetZ0QBf
WUI/GTbzWaYBhrD3z3KBJ5/aX4IXaKLyRRoB1+5fMBqHfHjOYInu0J7od7UW/EP39XF3zw5pKU9D
jMD0PiGSt7w+Hqh1ZxjQxw96zWmcyd5u9OaJksnMIa7iisw2VhGyAayqms824yOouTiC10SoD8mD
pToMlpEFxCwJSN+vdIU00tOWrVC0isMYoYGnrNUcmxeA+gBLamO710JuKpX7wNDHR0GNYJ/liQ4b
8UOXOCwrVwBYjDOMJ58tNSmugtkzHO5XTfVbfZUnHscClAw6qZ1uQFBFudUJqHodFVF+YfPtI4SF
LllZWF2wQOvTrv+Iv0OkRqAnDX2kOaDxZT4ei0Y28R4rJ7woPZN9KM7Qxa3N4IVBXVTGxfZowDZf
cAlltB6Fh3qvHzGk4or+K1lqvwTohf3hC/4eAS7pfWWuWLO6W3LDbrPBbpWFKjSYpwl7hUTHM3ZX
/HBGR8VmiosxeQIzgErgeBE+UQ7tQVCm+diCBoX8opglJKgV4F3ZUJNNteGTIUtNAEUU0S8eCU9W
u4sSj0EQulf031LBxTimEdabMww1TWCK4xLyclQveoEKNkwpXc622mZp9V5RSoRgbD9FDomeSuEP
tSl2y0fQ5rsaZl2fmGghQtOJVti/gFLWyHKeoZOsdRSFppt/3o5YHLhOY1KOEINaqxKfDwz0bBld
RLEbdhEw6NkvAg+m+y1+94lcut/39srREBGRHY+dgh50FweWNjVLlub6TcQPC9BBdNFCiO+y1kH0
XxDk8Ie4kUNUMIEuqQkPMizKwJ+KjQeux4KNBe++jcMlidrmlAbjp1DgL3gba7MWWgX+jPIfMdfc
ps/u1cNc1I5dsJUsMJmLaFiz7H0OC+fUhQe6xPniwjpQ1j9/UiCPehV5+X07lQWAn9gK7GDCe+7Z
sG35zmI3JCOCVim7rRPibGXrrYOr7iwUV3iVH8QIupzEwgvvQGq8nV+v3fNwwo+Ma04HhOM+QQTK
jmead0vrhoS/k/8PbRc4xchZ+DOeqqXyYs5t5/0zn/Rx3fXWnoHA+8yoR4L0FFBq8gGoIRiCCJY9
dp1DuY71zsOpLIu/8yPS+9qpflZnced1opVwGDz7ZzPui7iG6dEb9ifLgZJ3yE4ElV2lJZo4L7uJ
QS1w8Rd7giPM6B0HRokPsAD4SSPv1kBdjZ66nCI2OVMjX4NjJxHkV73SLSHgkC5oPVFD8dBeryE1
Ja8gJyuNdLEq0CtIo5Gjc4WkryJRVDuxBz4ND1TzzSsWwDD9OPsdt0o3BFHA3pb0OV+XXL+nhFbm
8ObaVnwmn/gQ9GglTHPYgAVL/N/apXt2b5XBssrgj9DqDTwrsjPusy+7ZCIoCZRbt+sELkDulY1Y
cU5M/SnS4wZQtcd+llmzlqYfpMkYZfF091jj7mqUwBJo6Wyw29rJAmNRptOYF8M7UFSFXPvbsRI6
dLEiGnryt8fxl5F1qCMeA0LV9ZuF+Z86kKoVo9rL7O/Cbsv0zNurIRLnWzb99mDmtwk2niFkGzc4
FlXxYD30CHLX+n9MxmgHt71CSwTMEyKtxp2tqrO576dySdCWzqP3SyF8RA5zIHYkI1M8Pl7X1mEl
5iilZxRLzRgxMpx+fjTgK2C6I385EEjXdxSt2PynEGZm1yDZFlAQKDPv3QUrK570LdXZPhl/CYdt
v6OmnbLiKMhbOk+6p9aI6RkLi9xvK0n+i+JKd3/vbJrf2s8umTF0QuzpomN/YveA6Tx5jWHSqQqq
66LKt4k8w5d3coUgf/p44P8Q8lWDWG4RPH9/DdGzxK5KX3VmqS4DQYK7gK9BJukjewvMXLpONiod
EaFrEbHefv6uZomozolwb9ecr4U4S+exdOR/b2PUTil+iPtlXI4RLDf608g6jBiZoA+LApPBCQsC
qBkbCStjRQmV8XmvR2jbGwsfkmxRmlqgQ8Boog5vNtfZVI1b0rUGinFn39qMmFhJrEjAmApfhHVE
Beqfgn+8ee1gsTnacL88cGEYp4WqGp33nC/lfvpIl+5Kxj2XBZlOfQ3EhyhQi0AvIIHMEHdNd9y2
NtVyw02If+aN3TpqdTuLpxD01iyrjTnfeAHUYux0H0KGp2rKLJMWDHIJVOxma9zQbUpeGg2E7BC8
xmDW4y4/MYuF++V2B6mLH6Fw7Fe5MGFreZipdGi4nHVKJKpwtmSWQsdT1eGO/PxLEA59rsNh/jFt
/IhWYsaZVQuW4vn52rdpzZnSAsDZ5DXZNOmBPleqGuwElYo7uHAy9vJTd+cqwlU5uEwOVnl9SwmN
uQZDKs5WmSH2Kxxvhk1I2GxcV5+AbYwu1Whlw+opgQwwNmlOTOmpHC6zjoavs2YZKxC6039r1Hy1
TtjP0O/ABf7OYCExqqUGjOjtRK+q93Z46P8kRrOgLLtslwP2Qp/KBue5OXgVKfq3SGRxIObtRUeA
ZXYmodIkCVLkydxrdZVGB2ysDPIUH00QdS7iHMoFBEc8LKXCeaVdLJT/0K7fqVSXs7AmuOl0Qyf9
z06SDh3K5lyBpSt/XZ4vORcXrEnWRPMMA6UcpXp9NGMoYxQBsvoIDd9Cc+QmCwRt2wj633e05b0P
w8DqApMiNSN/RB8Dw2gRr30ZRbhbTZq979AtLo8jPL70TkBUKVHsnfsuDlTgtZ2ThcbF+ZJeYKe1
CS/wKnAQJFlaJEflPuGQljEWmJDaM/oqcjWCN9tALD/Lpnz69i6sEJkoNe+b1zgJmp6C3CaMnFYX
93hDme2lK3O4s2kUrQEZvLowv+8R9sTvyCl5KQTQCCVNfK5+O1eY1XUG4ZjIwludzK9xYwQkTR40
CcDdrqCmDV7E0RixHOpZkZJqQIDLRNL0EA33kBgU2tFZ8PJTDgR4I14BjFfTKcu1euZzcO8Kdnh3
r+56wqhHHjLsp0H1+vRhgLMOOJgBAWl/vTZndEqsko4Cl5gln39YU1ySFUXkKoHax6nHqBIACmVR
EbMfC5jYnXH6assOpKgtMcfwHUtwx29//IpHZM+nMINLIDqwpgjn7dzXXCYZx3qobMN0yJ2Igw6n
AAbsTlNwfXi7V3Hhn/rPm+2gKDjlohAbhktdvcDsnI1s8LO0CiFaDbZhlR5XdU8NAK3F7mvPzpLK
/4Z9lHFL1alrhw8JWrcDHa+tQZXtM0xZNQlUpB97U/cQV6dblIYQVuHguZ2/Rh6kACUZB120VNV1
UCVtoaMLptUZKt/NzeE/lXA5dCX/w+CKc2t/XO+AXJmcNwaWDojNAhT8Htqm8eYFk88y61H5TeZe
MwEDTdGhswugjFbqF0eRXbT0MRBKp3GUvCuvfCrSVL4bjSYigpKZfmlWYSev2q8GsGialz53sQ13
e6fWncCkUUpBixWTa6ndFNyOGVVEV8oyVVHUeQ6D+weE1LuamnousdYNsEbnruiuOuJkYZhHKQDx
R1OCckoc+mP1qJn+hl7P3evkbA6Ezx3OVFc6GnMGFpqkH16hj/RkW1JUxeBhiMkMEAkAoOP2QbvZ
wYWG//gXe1/0uufGKA+SFHhnuLjl2bzi8iGAXRlMW6Kk/ojHKrX8+kh14zgwPOIX8iDO4aj2kM9r
zJN5hCxddqh/2N9tYst7hmLsvjp/MlfEktLN/gIOa6+G91NrjxY+AAPFi6GtxDNwD1Nf0V1WD6y4
2TmLdiINCJHitd9mEK64wJ6bQDH21b3jVc1U9DMpqXneHZGxwRI91INmsiISLDbQ8scTbHzz5mOn
7JdPvh6enkHSJv9SM4GxSgFpMapbNOoPiceG3gJWjV11udU/dM4ldvjGjEnoKsm+iP2fvMVzc+LY
nufOzSfeDiiwx12oQU0pDG6cMb8EPbtPQL3bK+CxybZuAiOqs/GI3AhcVgdfRha6QL1AjsHXImGO
70bditaaVYtSU6Vpz1CEqf+cqk3Qo5fPt72NWhwI3HIcCdppwvR7Hn9PibgN1yKBQKRocG5Qd5xe
SXEk7zkBRxOpyZ6X7DSTW5VQKLI1bbQZUZZTIJoUqZYBv09abLbgloTSLsZFqjAtgBCJz43kJOMx
jR1NV2B9fOaz8U54qmvQb8aq2f0E0sudVhnBfPABQUV/LW0lE6o4NkZMz+fYiNKyCGTd9aZqjCQi
dOw1QNqoIm80ob2/IFq9+sEA9AkYplKVdua74reucKrdEP7LhRIF/pDTmJr6MgPSTt6bNtEaNfC+
ViQC464hNkqkOuQzAmuNq0SqqyG3po5OBKCIMTLBqEmGuRmWCXaP5jT1QuXX6focNaGRVH0fHL3v
xT4ewjIv2SL5G6LtEOkvlOnClX/Fz7CV4SHHdxPDNxzdnq2JZCNsJ4BpHM2OhzJ2lmhoAF5w213p
U+g0IIVP0q4K6M2tvn9ydH2CB45aeUauYUuDh2F253w+BxL1nDkhqxEAGWpLhPOkBTAw1Gf+TDRZ
AM9fMfinhpVc4jR1a7Yq9FRfgpMMF89/7akc20FQBMgGa0vQB9ZYfGteQlbC8eItyxzcqZakTA8+
LKGZsQ+hBM4sFPsfSskuubJdD4L9MaaoPaJZf0JiCMng5bVy7dScJs0bPCc5Dtlx2gMherBs0ZCt
XTIIs6grkI7gLB6uPnu6wE7xwfpz3Z7eJo9skrSCNDKGZVpti5aiREm49xytw1H/yuDr9rDE/4Xh
MihClljoFWPThl20lOosBW+nPakOTQErA02rAxY5oAGXyjsddwMWj+EemNn0a3duONv6STrCiobe
n7hjJwd4pDZAKffUZiyi6/rRNqg2C7FCQ3RUiPVv3gSIfa2+cyBoiw0Cun7h5Xw7pYysas3dYTuv
Bf2nILpkRF0cNzDHxEIuKOFxp9dIIOczoI6sRZEib9Ucte6QXlgJo6jbOC7zPz7m7fPNXnm+Urny
MiOJunZ5mjcxHaJMvN89VBmtYU4z8EvH/9YV/qA/ZRN48O7/2X9TBpsFVMbn8i4yvyNaVQNgbXbf
616fW5JA4VqNz0hZtqpaZtyi1imraCMdWTwVb9YZslbhIuP+V4dxUhur+O4cDZvpL3UPwaIApqR3
jcRt6f6hLaZf1EmRbx+57YsYX5hHgHpO+ZpbOnTQLiQ2P2HZZBSaFwDyPhZ4KGvkqEqi7CpYe/Q6
qQtnuNwTvuOfZbgi66Sp1j0o8gSwFMGdrGnjev+gMi7K+O/1e0fNiMbdC/ArXvkRcYan3S4i8DYz
suzYGlESEOaGo7TnTWjsnEMz8SyRimjQAKIa+mNl6rPWTJiUdLKLYF/oJJpYhxQ6oiGq9YUDFANE
PVjJgV/qb3wwkMpJrg7bzfOs/G1/vd5EHn4FpdZ7pyGtecldinOhdlO3SwR+V4A9erOkDAi6xVBu
VjZjPUj4dNd0CYkDsglV0BajpWWYu3b/6JwBEu7nyMWDhE4/0zVWKetHmEkuB4sBgtqdx4Sz7kmC
jpLvMEcbXdw+hGbXtKjOOmXuMxatSumeAJP3d68my3qnsNawzngCLwlVG8FsqvCj+CtQ8APr57rY
NWSJhp0q8rs3hemDyhM2UDQb0/w2zpP69VLtZRQLvCfkfyYjrPFGlAGaxtnlAUMlch++0ozcxaCo
fe5eAQ5ERlp+bbG/vfe6V6u2GYC6nNuJPMdFX7UOE6/ny4KcF1m+BCRp6n3K53QhzqyKSSnv7+Uw
B4/u3zwkej4R7rme1Jvm+Tt/pqMdyzeyeO3p0yn2KyHJxHoIjc7ygbLrclux8ftpzqq79mh0u6im
7Z9VQqywSd/h5HUilN+KjM//tBBauLgmUd14uEBTMJcyWhBX3JKos64J7bsgFm6yuQ9pjdxNNbEG
eL7xqtURAOQsi0Jbvl/qpG25BrhD6pT9r8u29t3xTID5CGNJZkSjBIwkw2D3pRxVMYcTOMq5DWQ8
7H/mUAluT/7mTUkIy3y2IVT5Q/7AULE/cPrMNeAygLWFBbtJ+2OGRNjmps1oCS7niFkSKb3AJrKf
UyYPryNQRcAANZfVN067qYJ7Bt+h+XKHuRstzIk7IssH/LF4B8AXklNxB7E56EfdtswOhdgVcxyZ
WZwLF6+aiXbrH013DixZXxaKeETKuvAYq/3P48zG6mtGOQXni1era3mGkyB4VJ3vqnPaGy1JJ5hq
Ww65DOfj4lA7r/sJIr1K4jIY36eGXgyrXLeXMYfVx+dCgOsW9iEcl1P80zLF+uIgKj0qaqFYto5D
kGalgLIhCe3h0Ii+q+CHjSk+WIkX8RA9OGbOhGI9Hx2vpuo+NMBQ+QDIE7M6WxuS6TUor3f9NYxC
ish4ud6wzytsn5s583SOgN3LkKeM31G0KYrbgUsb1K7k8pPemoAhTshqZtMFdwNjjB8QMCTkuBOe
cKV9MC+yA37llJpnzxX9TJud4a7lwHEwBZfyWhNo3fmayeNTJV7HtBvHarHvPKmQpX1Ofir85mEG
tYCqAGgM6IecIC9GN3TxilOpCe+HFubOlmLKNf05rvoA0lCkzqEMiJfa6JN18byOasgSgpGDJfkb
YmoWNkU5mlukE6owTwi3poOKYr356Zk5Y/uDZGcpsF6QaWH86LG/+lvLV4OtV8PaUcfrYr8Qd98e
PdRZ5xsVAcWHhMgOKhIqlSDp6twRiSWC8FqBKQHO2YfdyJsSl1rw4drmGUgfJOF2X2mJZgj885v2
15nvpipL9/uIqMwC+ppoQ1T09hV8sNZIL/RPcQfaTwguvm+JPb5HSKAXZWIV/Kuwt61qQujXPUql
sXdq6hJeWI4CAMbtTLruNJkoTKMYeWOmLH2Zo/aBNvjyFlcRVrw5iTy0UE2r3GhxS0gi2icx+mND
EThOPGiiJc9GlXzr7L0Rb0dNXmv/7qVJfJc8T+NrAwZT9EVyx8XLrMmWX4lJxENVBhh7rTBLBBkQ
1TPqQ9mBRuLUO/v79OaN6YZtzlrdVPM93t/uQkl0aQ0br4mISwvdD9/GUd15g9EMPmbm2jSaukGF
bYkrHGLsxDGOhwYqYeMsbe4MpbPaJMoQH2ReV7RdSMTEYIODqLS+P7LqDQ8yyQIFYRjFTjCxRr1x
cU+MiOBH8oAkclGZhpbVVhfF67DGC8G07vghRsjxoZFXGYmEHEUYSM9htKTwczeBLJMUcUI4HFaE
jsH13F1hpnNJUOZh/Kz3RrorxOR9h+83HPZxGTzRNofnz3c2WQi0AIF+v2283S3Y42Ja08Iq1/sQ
OpB0EYZWdmjaRV7dlqw6WgGBXwJLmjulDJdp+Zt4/QGxRxqVyQn5im06DVpW/39HOFNwsBy33vEo
zZ00n5YDsCsnUdwolPP4pN/F5eOllYzFz8k5vplyByiIExIGRe5y2xEOwGtFChMt6vB3zwyiN/FV
vMiXQE77N1EVKyL4XfWRtiB/EhV9sivczJF9ey+/rBjH9tPpgutGYiYHsMy7+gOPIqQkYCbQqmem
ZOlytqLleiz3jnii12DaE8jtZtM/3GB0KEE5unu37BxYvOCtTUY/hGDPg+MgApUmLZ0zsqWwtlkL
AjxH+tKsIFOQyh9hk1SoipNbvdnr5o6Q8ZVgoKKuSMKpEGBqO2mMc7rwHsgXpfj+yqBdXoL5OY6g
/JerJfS6yCiNWCQphCbrM7gtmyidyI+kq2iWfty6USy+jTFkcBrhZYBsX3zM2DlJbgNFWKLZVGsy
F22YEV9dGIF85Yw72LKJ5Y6M4otokQlEsmEccyA03Sk2TkZf7fWjVxOsyFFSPS+FsVRWFpd3A50H
FDlDtCH/R8eCZZt+fus1SHLkAKkF2nyJMYkLUkd2fz7S4UY3IFFH3uksMRq/RcuYShtNgnrdvlTw
wdRFNliAAMuqSosK74O6h3DHnVbokSgaZEWcqxI6KCOzFEAFz5usOGsxav3SaPb3VXjzYi18A21e
GJtdQ/OpzSX/99Z0INj2fsTPMRf8/BCmrTz2eRd4Gi7CIpLGNnuNeYpIncqfQf1x3j5F5JU9mVH3
VS3Sb79J2743yM36RimCeqOzJ3ErMYVNY/UstOiAfffhdPs4SkIxNFWttYLEnrwvcolY6fTNbtTk
viId71kIx/orZ/Y9e7WdyzU49gE9IO2ILftw5etHQqs9EFgTVmHd/d/hthRIG0Dzs0uEFKQRpCZI
v5ynPAMbeeTNk7vX/y7nKivDPul3d/S2HsstN3rqMYodmQnnyBJF425m2uX8zd7qOT0T457fIU4M
vyasHzLiz3mS34B7OH4bTGQalmZqyhrcVCh9lxGexQiMwUq9Lg03Piw1NmFBTU4j81NnrTgem06G
riM0pSOGTcZuvUVTInK7ExXp/yoGZsMX352LXzRTWh+Jwah0jGKE08/bGBlo3Tpc8cJgs/g4EHBt
yWDvdGt4HfyanEPeCfQyNJrtIWbMkln4Ra11/4IZNGKVfGiOF1AZBHEf7ceVScZzyCMtBwWx3eNw
tlU9c67dAz9SOWid1wdWffxB7yY75jQok5XeW/uxMtPysaQmGpJxNnYMTEJuGy14BFuFWQgm6KEj
SNNREcez5GdY37nqJ6ktQi7XqELZCrGAXEGP2Js8/0ydCYXgcqm0ksJKz+jgUQFnWIXPpofSv1Qq
u1iHeUBzDdBe4skpWBUwNy7fdKEx/gngi6MkJ2Jn8AEGApQgr4qUdPpU1KPiYXs71aYBmRv7lKe4
ngHsbEwYK3olqgcnl+VvFpftfpBs6znQ3ITNP2yyf0ZDM90639wezBt08YEhk6GUBlsflwXviAyd
BDGBNkG8OSfuhR5KcBYZbopz9pBTG4soGY784q21NQM8S7ZGvvFofGUJqdj1Ma36cWuly4JI1Wtb
iaPIkeL8w3urx42rrQzEXIi5febAOAyZcJuZikAgacAOBIkmUyIqQcYGh1EZbR071a/ovBHp6zIU
A4tAosYLUwWFQI71x3+PoS58QaY8svu1FAg7YX0dwmye7XNBC76GQauAbBiBdQfMmdl6r/cPZYBg
VMknwXnNy4a3m6iBYjcD9JNdkw3bALk3noaMfvxObfjq65hkIUoLpIQ2157TKKowc9XHzylS40nd
7qmO/zgULYflyMvYnMiU2uQfe+ENHoCxn4foZTMGJZxgb4qE9rJMq2TY0hM+NRL17CtOMfDRD/Qj
/J7VJp5+Vc1L1Fa+YjBPU1UiQ9XLBSjTnB6+J/QVvDPUDjig+cIZpzLDvsN3M5dPobIiQXz/X5D2
RTMQjnbNvR9m2hEOYqp8NNgSKuo/T3y1IUl2xk/XsLLIXI2obokYJQsK77CtHa+fMJ01FcW+xLTy
Sp7XbPerHs4j3CGxBRCXMMR2yxeo/QBPFMiDSiwH7B7P3Q2yP3MW4NiSYEDFRnaoBtfrznIK2xF4
20hvJ3VCFvhT+aziKlIee2xfzXj7ZeDrhNER+D08eoK3b9FkIIrY1Y6zpTD5Gy85BQHN/rIpSS06
Aw/nWA/Qy1A3ZvJgb/oUpM64ymSdHJSqn0agQaUjPpR+gbM8CLMij2PYVzw92zl+AvGFrjU8XuBk
fTpKJIXr1wXFzPdysKOdFnxf4w5V4++9zfQeaSs9ENKarwUSxxrnW8tfLRRkZN4fDi3rUs6W+cQq
QRY+mt24px4nR5eJkqkVXYR4D0NGWRXmDuMwnBcK1+xQAusJqkjj4V9EnDgIlWXdTfJGyKN+S3LL
rhKACzmW2GNAgnA0c8qGvthoC6b77SHaI5Vp5h6cRbtS7I4ePv38DA5W9YxIf+GzWr37og9WhqtZ
pTCiJu4Hw3AYq4qEW0dazQ9lVoyT7Ug79C6n5Wjh1GOhqlL+JOS+oXrfr+z5SVl6nc3tsi4/KkNd
iOXMZnU+8jgRfA54jjUhjb10+W6rF6NKPFUIgsbKnLWmZTi5pzIOM1HOP2T5O2dkf6rh1YvvYN5l
EzR1bpVebDiiISsoBms+XxNa4U/3xwOsoIELqzW4HhaKtesdzTyKFn2GQVkjrVKZS+L2H0Dz0G4h
cwO67pBXDfex58OGABoOEknsHHgWPRn4TfrLLrrDSWk73kdLUgSYA5sso3/ECkegr0YVD2T63xvu
zJsT3wFYeaVQg6zUuddlOneRIu2nWnQpuRjSoie0VZdQ6IfOzLRKOd5iKfcWu6okPzeB4QrUF6Rg
6hPtCdcjlrqnGbnIQFkN0wEreUsNiJrspJEYgOxThIqyLPwnhxG8Tfso8tgGlEtRkanvUgaV5A4G
oGKF8jNXxTW6p+yb6N96lFzKQlY2/AR8/9/xFcD8qspGT6MHfx3hsL2bIAN46A0qk92K7qhKVubN
8sEItFeVEjFqvZV+0Lso/au+LLOnQ/uNOmIX+3K2MX3qbVqeL7Qp8GfV6NZSWYqCC2uvhVSeoZra
FW9MrYyiSYYP3F10PmDRJhn9sS+zzonKXyn7G6SXJOBihifQUOynVDZolWLru6b+/JlPDZa4NJzo
Aelrw9KsrKFDxisLhNUnge3pZzDlXabDui2OXknhkwKyiaBgc7EbkRRP0IjSuQC0srhSndPY1ERV
uylWDBoha1XypK/87ZC8EAxdcKIf+kEXzoLwVz5CF/CmOBBdJLEbm2MITaMSSc3Rtbl2yTnZhmbK
P4kWtlXvaG8odHZh05cYz0L0r53NPdTgWgNnRPdjSZ0EFSpoiJRLxqlMha1FwovMhd3mo2qIyUvN
zpozT2fzrpAwB3jo+yPkqj7r7eVbfI/M0KxLnvrz9uV5QPF7CkzR/iFLGLKS+dFrbZX3b1Zh7QqJ
Kh07opZBr83h6muwwZ/u/w95lrjfouydmxOK1abjIvKgXEGVr8wOKD6lToHVklmpJVssqKm6hh/Z
VAZYHzFq8ATSE+dd9tzYvRac7NhIy5yOi/q+1ni9BnHuZ70EChwaPTtFzHAXCHvyotijf+Spotf2
6OzgK8gxmjyh1CTRFC923sN33brGPp6bR1qQNC2tHa6G11KVw46MoC+4l50jve6egq7v7JI6ClXv
jgVoM+P8FeWC0Hb7qsDfctY30Ffko2TFqdHp8FB2T18HI2faad/OChLs/FTFcPYNjrI3V/otlgHI
eZfIfRTDNtB3dkFJNeHghvoLWtSD3QQOh6H/ACcDbjygCVgsp7iSSA185hTCv6UU/ggqtnXIVR9m
js6RJBx2TvWdaPGTFpkOyYaZNUFtCYHuqjCLeLH1SJRCC1sLe0NYgVCtayhKAXYISOdpI9hAAMme
gWIsOyEYM1xbw/xMr1z7HjkK+Nigte8DNW9TTJo9Kla4H+NxQpYazDCvDPnchbPlBF3pfXlZ2WBK
WoceL2F8f2wlix4mZ79XQyu9kRLZ8LTGVWsUotAcoG5LfVZ6woUkHHp42AAPlhwAhmD9ZIkXdmkS
VMXXoc/LAevpjpGtPv8DiUZKVDLByfRtHh9UcRpT17FjzJtvg9Qgu6Tt2kkYBXFDaXZ+XkYjzyxR
NnILdYAQTV16DHWuc0sYfEWGvpZ7L7a/y/ZQ9rbukmEz0vHp5IclbH7r1+CSB1Il1+aOqOnCa9Av
Uz1tfEgYwlqfC+7ptMb741rg6DUkT7DbcS6EdSl3UUVERamTp/IaSPQ8Pg6HBH6Yzxpvc7+oloag
AKIwBxtLLnHwufHkGPsRsD3rm8Basdc3LWvr01X8b1FJSVzEKQhPSCje9coj7Zv32R1WaBlUq1v6
w3lF4aulNsbPIJRlr7BAoqJSDl24CbVyXCpFKhA0Pi2cMlc1gQyIEQJqVGWYDjuOa+x238mpenqG
sbx0RnBOfSb6QW5myvGOp2PbuNm6KgnxD+zyKXBwEdIJp6MQVgY3Khhe4rw6AEJ/MDMmFpYjmLY9
ExZ1W6NFeKOZaQLBVKVFWFldY3IaSq7HPYaSf+SeViCbvxkT+firqTKuuHoAIRfC9j8ZYUPCcniH
8zxI5ownHKFJxsk2kC1Le63uYesHwBTfLZ3DGntpn38wK5FJ3BwBz8e7nGabmBQ4Mvtl8VYtmEsV
8WiK2mPK+rkeJDJ0EsDizUZyagsbahNyKc2wabKJX26+x/VGrCXtDBPBeYkQFRvg19prNgvfhP2B
VgbDkUga/anHRaB1WNBopHBWXdJyleQFsjn43QaYHtce9rFO50VrcbCYm7VYJoJIsQUNzdCrWr1B
UsEpRyhBlZqnEKlOhVZZbsOHLz2+sFpyR4tJWK07Q8a7Yt0RV4sDrHj2aKZw5CPeqd8rrefwMbsK
AlxrF1lgN3hQd9vZtDlxaeCsvX7VSNIH8l1p6+GGRAnlY6ESQrVXUufPseF16yhEDGJz+RjZ26dp
d3TwLD8SF1rmjYMcHGKxiFri/+sA22hpvqBoNBm3aOxo7ekRO4SERF3bL4BLlypnBMHikYJVytIV
VGGypsTto4myv6HI9E3MDZF/RYLZB7VgOYs3knosTcf7Yz32GO4PqcX5XAokWEPeDgcvk12CXdg0
ulOAYd9GrtBH8nctD3NpwzXC/r86Mqt6i0/XoXC6mRItVoe5lrE74FNKVeQw2eFYkxOPlMJlCXyL
c3ZR/q9BQmMDnG+YVxGa5AD6vTeFBluqKHTJQ/6ciVTv1uJOlunGxSu0sIH7s7chFOAZOTKa4m81
VGK9DLlSdnAt7WbZDYq9gvlsofTeVcosXI+8Dy7FHW7NJWAnLwIK+WkrcXQKZoACoBcffuNl7fsO
O3ItAFVk7lXQuFKVXWPWnhBUQurjoxz2p/ibDHH8CtRrUG6FkRGw22xevORjK5Ry/f54zut0sYKK
y2chTnF0mrxn6+GMLe4QWbu6HArziBwIUpgs9jvnlJuMTOpBvCS8K5rSoDCKoTyAAr2KR3klxNLJ
AcSIJvrWnNZ+KN/A8Oz/HnrgRN6BkWhqHQ59u1K4xvKnpD0hEm/XrYXlSm0NV/Xnwcm3xCCeHa23
h1EWq9zln1a2wGzSuIpg8kNxMpUUThLkneLhGGQzTn4MrCNp1ET5VAlJohxPC9/mDW0tWLuiqsW3
+cfSzdRVLbOYvwXrL0Mbeq/v87FpcncKiCuQ2XWc5mUEeda8xUJD1KDqHXF+qdcFfCiL0rE8xAmZ
DIts96YZ5+ByNfLf/a7FMXkJV6X2lgKzm5PAudSzA3bTEtRugJybZVnky2U4BnlhLSKCJQ7G9JH6
BA7C3gB+j6PWnLxIPWYPTWfmuKKXystnvHtmA1GZbztvtKf/rLXQX93vqp1zBwEvh9cUiUvyO5pD
IjMSXJbf10L2Fbwhd8iVlZCFgTVeSa4sCrje+7GFlANrX/drJo1Uxvbf4Av7BQ0UQskR/AWRH2w/
6PhLGaXnADFqt2L2FehY8taFS2Z8bttEdFsm81NA2GfTgwaAIXZozZkTdfYaDp+fz6u6YCQWreFN
efA3jwJtYEJO3857XIB9jKC55nAHKEE9n6gsT3Ke/etdtA+NpMhlc5+ei8JHvls2EaI4JePn6jTQ
ba4iJ0UDitvDRPcurllEibDXrrN5UlqiszyPQaJcI20YqSQIZh2CNYbqz+7ssotJfen/8rwADYPK
BIZZN1DoAPMi9BDfiJMQhdcv1j4o5WeWWIoOtqSzd+urXEPenlDKFCFX9JoKUMtExVA2IL2neMVe
xPVb3y0O+gT7skJ8imBFy70ioCPjwMIuxGYsLJv+Z9kEFSaDwRfdyhcW6iYlOYReX5aum5loWjqn
8nnf9As/3x4KzWMooeJ/trTZUHOPocG4jKSdWYTF4MjbA/LoycQgxibT7fW8SsuCgJJ0LB8Vq4sI
Rz1TZAUzRtlmYrzHpqGe06mWZbxov++BvF+WAiOLV0snlKVu97T/hYMNnQ7TwYFhWaIhKXGV23bR
zKf/feJiWzd9+1iHSXaDJc2XY4GPbl9icSR+UDcUjKUfDY1hN711vwlRNrIHRU+lUgoLkLiHwXcZ
jb+3b9IvGbMJa+xZE9b7RVC/v0qM6IKBT6zYbdIaFv2u72+OmFesLI6xziA8wQZr2alZv5zboOQT
AD3z2j0HY13jCb81ECyR2xhwfMMRts3WCIPm4DInvxPXcE41+LP3cooZ+UULAb+YpcV2J95q8YB9
u9dAv+0XPzL70LVpXUsqHV58OGVI2HAubQE58kzdG9/tzunXW0L2trH6t5uA2u7GjPGSxrUmd1zX
5OJrkHmgA5E+t5ZWykdDTw/41YogeGr6nfeJGjEImeSjMibx8rLl/LepSBa/ZWwy3gB115Ot4ZI3
0n/jNrV2T+kXBSONpijaNcM6sv/gyX8MWphyTcTWMsQ7tq1i8nGF7/vKq5t47K37FaOWUNcnEKR5
1rVM/BmiB3aj6b4wlKWKuTfPBhw9/fkpJITM9mGwaaO4vPcIIwvQyB4skAQ7syOgYJyF4uNwFmmn
29Lg77nGBcqrVa559eeB8md7VqyChLXtkC7kQSMshQ9Gd4SCnQhsniQEdd1AeVkoPUqW58YRkfnN
kTlNe6wULro8mE57JBQSxwLKbc1NWG14SpqQxX852n/LinNFk0w747akNAgOu+xvOd+volGN0Ecc
hTU318tgwgvPH/s2OnZIXO3yP/vJoPqPTSD+N1C+UmpyDyxEkDuVVXXgxz1DPrkR5q2eBCQJZa9Z
UMEMSi+SwOiWpO3NKwCafyblo1q9XdrnKMtytbNjRqbn/xritNN8a4eFTeM8qJcFWbDjcP6nWNNd
v112F0jPRDsQXhkzsmCXoEexLjvi6wGbUoOL4enKMixGz++TQ77eszCD3Z/RyA9hZp4xgIXqhnkv
qwLLxN9D8uJIpdAT0ZvBp3SV6oowpZ3khC+FdgnTNK/5Y5QMMCIor1kIxmZW8zNXgqdts+bKpN6M
+8x6jLV5nrN4UgNZ8eZ+IotL9GEjROmRJah5o62hdDqHZTEm0nN1fO93inbrsSnlA+e56dmh6JZe
zNIQgdN1BzMVZfefHDUz0FZAWC2UBrkO7ORvV1OSwWVjoc4PpOjdiMZA226jOrk6yX2myvH4PROh
0C1pbHiJy760cDKajhDe0Y1p3p+neO2gZC0U6JE7mDj2HCEmNzIeiGrbxFReXbs9/e1JZN48uqx5
25gNGcctzU6k0lm0CEUqkmJT/qm0Sg7p7z7Y5oIdmJysMglJVQPNIMZ9l/QTAMUDrSsUbWy9p/YW
vBa0Cr1XXFD1FLvpnLu1A9NVtlPZ9I6+p5QtxvlzjSq+00CqbhBFKgwMXu6l4WcDuQjdkxRrlRnG
l/0ccSDIDgSVFucVqtex/LCmTp1lCI+LfPW55RdxHStRgZ4tBohhUSzZt5ZkmRQ5+9K0BroZA6kV
kXfwc/g1WEX12/37iZKGD54s5bzeWqlkIAfTz5DCf6K3ou9fclrDe5I0O3p91+Y6S4gxtW9+xH47
xQUDqbW1fcBRzzm560Laf5ELficeYv8VvOdiOBsFtngbThbHrpT/Sseq0ciC0rx397QwdKg/Q7Va
XksW97NxGll3tmYGTIxU24CVd0T7CFGN5OkzW2jBYpMLqZUGUFuq89cY+fnb7NyCRBUV9Nm5CTVm
IBdy5aVHBReUYTZw9wfV0fzzJz1FJvfbEnM1O8E1hMKIF7EwXN/JbCcsfj7ZY9EJv5djtgtOIUvv
AoNiiwA4Yp8YkIzz1s/Y5aIFCUK+LLfVgOZFl1NMpLu/71n13zQjQffslIO/aZY1ek7MhnxXIcjx
4GVEojTaEaFfdbBCJ1yqGL7X+8veXUODULTGqhaQfcbHW/O+C3AoOvPejQpRAMwvDtr3nbEemkwV
hvXbRb4FztS8bFo+OOFR4Nhvpen5bzM4nd+HSoZRTsHGdKm20yCQixEATEEi6SO6d1q1GPKbD5sU
czkqWLyCRVjbV2YmBwAlP+OpxyYz8YPHmXcMRpyRffUHiBMBkvDeUoSewDL9os7TY6W9pefSP52i
94SSOv8phEakrPBgcCr/KelIspOrUVsbGLlzzfGmVPKVjoBCEcpds+zeBQaHxi739TIaA8m/tTBX
K/4TsIYmw/kMy+21jEwkP3XL31sbhucAj+O+4sGURdX/T5eORJTXFf+lkrm+m5sdpOWPkWf6NzGj
qyr6JmQsUSR3o29WCyOd6j/YphSDrQvGIBVl5Gw0efBmgIFELU61gqGw+AJfAoXg+vtLhHz1MDiC
eHG+0XO/vSq//xWfznU03uOQ49Etf08sZ2fscnToxUPIfI0IPdBX9AiQ6kdX3b4UjK4SNGUIzpEP
f9i6Z8y7bgNOHoSyEpzA21bKwhMRm/6vGL905QxQrSU2viAYhgBff/pIHYk2DUH+UgkfzaCTCfX7
PLOgmvZXohXpwVD48enoV2i/d1HCzWvjYAdgDdB1ocSpRMrqw8bwyhiolGWk8YpCCg+NLzLWc2+J
TmvaNBP4FBSiDRm/T+/DQvoyozQsNF1f/7pb8fsJnnGEcBqdZ1p1xyxioQVZBVeu2ScHqqUUM9JK
GM/eOC7WxKQIufBnSvfTyIe0zANAiqKA6s6qTamsiEh/oiM9B0BRvBk3yc2WO0t53aw7llKAZFvT
YnHv1adsuc8InyHKQ7LrIZrgUWAB0DoVV+dIKvmc9ZPyLxzYUfgOhuKx3ygXPNNnY+4fKUlD6yeB
/un+4xNBNSMQ4eVVESvIccTB8TG3+3xXZ3VISGc7NYigh2PCsbIVB+OcPKiFN1EAG776jzy3fxUJ
gUwrZ6j+oottSvEXGgzNPxrrn+2Ix8HmHNDLXBavn/Cpa7sw+Gp4kgr3BZoYlGWhMUsIqvAl5qop
FJ2shHXlzWd5YNiGT/DiSgVzQtUkxOAd8H+qr5Aa3j05FIM8rBGeAF2xJFoJzkNYEtJPm09de9ns
6DwG5C4LvhTcVPh32iL5gKxC9HncvoDHb7qX9yKIBhZqvY5WT5ANgiJ/hzQD69oVtsVzBF+m5Iuv
95d+O0UYYU0jXm+z6Mhz7J30L+txEOqF3rpF38vH5JRmPPehCZMlwDLK7Se4xJ1zh+1nyxVjxQvA
8yxGvbTEO2+3xmBarC67r7QZHPW0dOlChsp2XqCxiQgl3y8R31Nie81VX/KZHoDiW/J3w6zuQ9vg
NhjEQqWjkGrgwM7WN3+U+3cFe9cwW+ZBDZK5x78YM+O65FEMAZ+p7DvpO3/5MXT9LrzXGt9SevCx
kInlMCldVok82Wz1m2Nr0vRkjCZUDWJHKWeEAZ94/F+06y8QYemVx3TA3/uosWFWE1x9XmUwpe0T
6CeMhTpUzDMkFXXTUDkh+jebr9B7X166e6eMiKk2qrRCXOgd1kmgBVkt7TEK7ceQ/8KyM7ct+BSx
nC8ienlRNHe5W7mZQM7Z/N5YyXWOl9F4mMsz27q6fSylKTcMVe43B7A/apBqJeNxj9egbX9nXZMW
GuTox5zFu75xMb+bLoMDNGg4VYrMhQ3CgERmaT1zHcscsef+tqQv9cGt2IbO9p1ZQe+fzndW8DqY
HTLXW7YetjL357x4WeJxxD+m0reEawpRlmZKb7zb32QJm2FbJCtpPFCDkqrOx3LJgCDFNrTIaLZZ
4649XBhufHpYnGFCkiKXEQZB78T41WFEgYxPPhKipCfSabFH6FwP/3XXDXMkKWIrLcjA0MvtYw1Q
MiGBqFyJmQk3jl3oUiKNXQQ/9f+Ks43oQtFB45g2Y6Br/isWBen4j/84V6rSPgDQBlDVvLtx5FRX
Qim/CLKDdwxTW3+ibQcmtdlVBbcjOI4//yYYeASTepG7yKCNjBO95JJX2mr2Wg7TzdaW7BR4lAFj
VFLwpkskI9HH1CXYbwu7fTGlHPm77D1gF7jjYvuXmX8YgZa98Bc1AHzPX9soz11k3vX2RuAwthf+
axz+5acqTMZVxpARu3WfD5sKqPyfDiwkFHvViQFCuuqTBgR0L4rGN73ovAJ6FTQ6SY5s9IREIHnV
X3EngzIx2xfgZSunKaOZHUbg8OeXzCno8LdheGDQmA+WxNkuKd3rBQ3IIcDqqAs6pYRK9lYo3/s4
Mq1N3ucfctRwoSnIffUiLfCXJyzwcC/+J75NmFVb0N3jwEWCLL4sKaIvcWuJ2F7l4QkHJ1IP8EqQ
veIQLJNb9bVDu5nhhwosY4cmsctgaoWJj0wyaK06HfffY0GJ7UZiXs7n12Fki2hpCsN+aU65W4BA
rqcJjnxgfFbDchCNfUPMDzniq8kQOSPBx3zwFDyBiA+AlYIpbCdlWpfPeAI3bUsFLCzIHQWwmEa/
Yrxg82s7RQu4drI0LKTZLhpOsuS6Tv6fojmQEnOUsR+1pg+Xdtn2sgXTqEObf9FUksEveTaruCf6
Fjio4jrMW8PLHz9TGZ869dJUmk1isFrM+lMUuCJjH+N2iWyFq6MMRlfvhi/4v7nZ5ig6tAe5b8fF
mWGC4WSorQ5WuwqbJ478uYh6Q3NotgE7TYB/iS8ronwaqrNc5QlHJHASqS5QBUobUSWt2sgOvFwl
7FO2VXrycE/9gLgYAxV0HkmQBaq4fEFB0B2g1lDStzlgb0F+K4SEKbL2cKeQ4+ouw0G5SAx6vmYG
tRmn0af6QgxvyNIX9G0O89zgv5v7WCnBwiuH4EfbE2igMpSARnrTBfArhRg2F68fDh+OP9nuPeyH
QMYUrNtdWB6R7yKgXOhrZtzJnIGuLg44C6JYS0EATe/Yk+7dAMoYNK7VkAL/LuN469hCVi/W9bKT
RG7U2IqlsRRnq5gfsIfp1te/2/MfRP/w0OfVjI2whOgV/f9nTLhyBQFHlOiUQOLx1TjCDoHZZS2P
MNE7iV/jmZ0gk3+ot9Riy6x3phuOv/3/GJ0SoUpP4JgkPBFsiRFuxbGsDSznsvp62Pb4w4/4qDiX
OTPt92GYQ9b8kDM/Bg4CNuQYJjez6fqRVo58SrR8IM1mMo9kFksGTcdEhIByIOHY2B/+zPxEDsRB
O5MU+38I5zYPsrboFBU7MGhWj3cdOYr2WGObmDLl7c/8qeesJDy1WSL/90judkJAOVLzl8WX0FN3
YPT+mKo/Oqo6aAcMX/PhF2Wacjjl9NvUnxcvavSlPrwELMqHFUwORY37ruyQQDeXu4mDHRuPU5XP
IR9Ljl4xg2GBhD8DxwHmGLoM5wQIdhsMytyVqld3YD/MNQiDp2GkGpXlCrjza47uN8a3u47w94mM
G9LNHyVjHfViBrMfOV5sWJvw/qe9/oJeC8Of3b2JdMoJMVnLjw0PTv396qv9soGBUHf2SkQpgmZV
1R1hfpgznZNn/VyrIWcEc2MgTEPNmqPsQgosTr2weeG89ofPyCt1kKFQAJKrYeY2ZlolmMfRtq+P
cpihnqfW2sFetnzGYL67tg35ftO9lZO8pO4E+i+mQGyncCAX4Pkl1334smDnx1nbyQC3wUguRs+4
8ts1eH/hVthEuLrlm6pEkuLGU14dL+vx/ofGYwTXVFHxV2FBMmMx035f+ywUJAk6VgC7+XTGhw0/
pFNq8uiBuSMDrmKjSUVZgRcmavRCIzPZx869YrBPyPq9wsYLBs0i9B9TKmZ9Mrqr92DLJDG0Flmj
9BPbz4kPr2dxdNaz041mYAGfStOz2KaCSpy3HAc6RxSEplB+d3qPaJjAvp4ZfRE/XAxxFPyVp7FR
SsL51EUmuwxERdiyyWYELe6YCMsQPu54oEat/I8pTeC8tBz36WkuT4lhEw984Jv7v8M7NFEChIrm
iDblhigzmx9qP75aGEoOd87yoljmh9nSTVAe7TInY5sL0d/3E6XmwHiRBXkok6YHPDz9h5yIqqW7
jlyXBd077f9sXRUDlWrRXq2c0XOmzOZIUvfFKzAM5RrPzDHqEhhvr26W7WRMvpY+NTfyjYd9Wj1I
JVPs/KYuY6pAPjwEJKgVw/VYISEXicsRH1T1zOikOnzwjCnx0GE/q6/6EYlefYoezPNWmUlTTLbg
UrFmg2BFe29ShPfBbaLQuYdAncZSWEOvemohvX2LPmnyBUeI82KK/tb2NocoE24XqdwQ9MyEldO/
F7HslCXEwOcLt8WBXfPpL9yR0YTM2D9bcTWve6exuk6Fgc28ofGRps9OyEUQZ3quRIpKxKklHaAI
vqLfeGPXQTgI1E5GLSAKbolxTzO3ITfICXJ3+VgmiqJBEyhiNcjbNkoFKaBMcpQsnp/QjjbV7RUJ
MRWfgRWvy3F0Szf3KfPtoFOq8DrCytPXcuhnxum8GjBX8s6RLCA1YfOklUWuA32RpzqaRAMIQmDx
cFaIbcIq9n+anP9tdG7Oy3YNeApV0COM0cQv8nnyRCbinkIFZu1KSBCmZa6Fk1qlB7CRb9RPbe37
MNiiwCUgUDoAuFndQBlwFlXtY6w4N6/phWni0d41UAZPOHoUS+eF5E8m/UDf25brlNW5teyrw9tc
z2ddEExou9zfSfkSYAx66+2DDOnLR8oHN4k8ViU+aA4H5sq0ZnFlWj7ZL/cxJ5eBKv+Xg9mOhy5i
RzRZxXV7EBo5B/gT2H8Aq4A+IWXL4bvNlqU/3ED5EdAYID75WxZ5Yq/K751GxjZ/Tq7wjShA3GA5
rUAR+fxfQh1cA3lECZEYZTMyXy+qP+ySW4h0tzXh4gtTC42geuWQJRVyYfxDZ+mtClaCmry5JUAw
nymfBjEhvwXRLLhB5qQaq4LJhDxrsC6HUU6drkQhDDwoJNpCxU9b5O0FXIenTnXqFISD++8ronEj
5gwezXLktbIjDqa3eE5UIkMLHty6LXT/GRtApq33dFR8xsQ3mQbcdDwOKIDO/TLBqzTk/5w5nNmE
Hvg/YGSexjp0nOhZ4BXvje6ZYhOFC3O4zMYWwqjqOrCcBk5o/iaKkiXa1Er8dIhNM0kkXumKhEfk
MAJOpLBe48NIWnfMGWHuXmxEAeyw/SHDqIczJc/OJmXOFLQ1u+aaTIQ64xlTjy8FI5cdX2J3HWZj
H9f89LI9876fFiC2Kuo3qDfzm8n57bCVgxF2gI5MitNMGv0swckoXmasiwoxStq2YT+3QvNq8XWt
pYMA5ky4p3RLng8ZfqJi+26qMWchny+kL71whQ3cjI8TWVXRhQmMNSt1LO0+9TQxZasR3elh0Kyr
k60Sq8JI4s1HnuNiP4rb7KYxw3ffXge0YogDqeVMAoR7Pqb/0eACLWW2ghmmKjdrw2mf/SInrwjg
/kIGrwZoewWhL0DuyBEXAnFtPugfWJ7KILTZLUirTEAVUe6d/iG/DgLyaI6FySbAt7MGSxuDfleZ
7LUyT7FOLzP2USPVrGn6wGAjfIG9NkZI60VBuuCOihixpiJtU7MbYUZnzG3XtDip/9EXHwDvKDQl
fLy7C8BQwua4r/7rHd6H4ansNr1xEb6pNUrtLE8VcyIAq8b10/DzKC5A7r/nMdO4RtSkoD/zfKUQ
iHar1YlGWTp00MbXtpU3wxig+wyz7yR7Tl8TBtGayTQI3+yaBsSMQWIWuzF3mpweL2wmtml0n9Uv
81srNNE2+1lKBXAUs8dpyl4lp6x1hZZeSeIs6cfkV52btEhWSkRZCYV9MKlXko0p8UW+oWOg6jiV
D2UJoQq5rxM8sZ0vrolT9qYSBAI11q0xg9faon0jhkr5QD6j9vETxolH6dNBxXGR6unVPrKtnhQu
OVlclruJZIw78f/oBuMJqO/Rz0qmy81LmPHLurkkZsLX5bhZNA63/EvLoHrVG4va/Id0aJAMc/n6
TylHAi0uYNmuEUomwu+wZhnK7tGqn18BAps8tZBW3xKVXoV7Fr/RuVUSflpZag/nRJ9CaOBws5vV
sIq5MmwxR0I77vuvz0AEPlTtd7VQ26phTx0/SbudvVExuZ2eSr3NQAZhZBZRzbzcyZYkykpcDYO8
Q2C5oc0cLGWyZDb0cR1J9RcHcghnp7Q9V2T8FdACrOKHoOS1hR9+Odncy4eykX9GFPczh7XPYUrI
t2/jvHJ1U12x6Y10Oab+ppQe31obs9SBLCe/z+XkJJOTGV7edXbMoVvD4JFinjEVTxWZPfKwFgNi
MIci0ZH/tlfegzMEQsqhtDIk0lWsVbgEGoHuOGHV02vsZWDzI/ItIA5t1o5c++8iREK5SsAcrQp8
GCecup/oQbfHI1CHgd8R6OTM10ooKHfdp9cqA5N5CGKbckQkP5PmIuvf0X2AytzAIbTJf+ZLhyi8
NRCxiYPzndFtmMWApByeKyqm+hk7gvZ4jMmh86AkESn4Qe78vji5VTbuBBo2oCNs1urTGDh6AGMP
WDCdxB+1+eKQWc9THL7NW/X/r0n+3IORgSpBEeDM21pIw8lYWB3NuTGy+DnjE29u7qnLM6jjDwg0
35mJixzuVF0Nw047chipibqitsh9wrpHfNZcEk/iyG7dxXymZ9JkFMFeM3AFZPs/m5ggqQaGEAif
OMzzr0pr1O4pZlYnVz0XNRjK7aeFZB84f2xAkb8u0e6v6Z44TQFp+2VaecRE9sNicfEw1sfzzC1a
NgrcSiiYryrdbsytimv4WjCYiEyG22+6ueGImwb6/xhB2Mf5WQBeo2BTdcM/ndnmL3uWFp1w7qQF
IHhe2oMhj5uPqUXcnlc+fpiFhoA8Z4Zqtjrqf2WoKloNFIPBWvR3bcaDEHKXzQJbOi/YsS7FQ8CY
NQmmTS3Gz8kkVxT7gUkoV9A1Yo/vSvomnFFoxCoU+VyErziwW3lcUOGzllNDcWoo0rDVk1L8KiAj
J7NhgV4rNNTfuVWhf7DmJWiw35hqGHspkr/LK6MGzBG6LCsV2kykWDOXfFgaHRsw4U+eLHHqFWWI
Tdo1txjVrKXTLH5wQFzx5rD8jt991vSae3cZsZlHbQgOozgTxlZVbcASksycXH92SoV76J1UOa9s
CGdh6NO1tve8lFbIpXd3ZZuWTraTGWpWcxc7I8Hq4TsawMo3Q98+0vSEP3N/Wnk1eze3MgMcA8Tc
8uQC0JcHAfWWRIplmz1AZsKFW4SfXPd2RnmEIzy/dRC8OrvlbvJ6gAjUSppMgZFxkN8wGH9wTz9q
IJEbQkJmRGhn9FSym2k4eBoMlVFOjziD5/tyG2ls2GISTbhe1+3SQ3u5d/6izSX9qnABBk5PjfOt
nwlYx8NbiJNWcI9v1mMsWy0+ISINDjJmll13/QPoqbzZXBszlc5n8NsaBWGOWu3FzovjQA19dD7y
uoemjiZJQTAyror5aWuMGfSJfFT2AYlxcme0y43u/mxU1GQCi2eJTcKRglGJETYYeGHIUdGidTIs
A9CMAzFpggIk7BDE2YyvDEt/yJbKPuLaOlVER94YRPCc+CMb1hm5shqrYtge3vjedKIq/sMyoXSn
DKxs1v1RfQ7ZXmdqjWcKYDWHr8SRT+iV1CW/8kho+Dp3jg9mDBOpCQeSEiAWvTj5I3FEgWKpJC3y
8o68CsHM45PCcn4wirQm4HV+gYIlJGyl/qnFoCgZSKgGXM/4G0FykGhAVn1wt2ICk10vHSvP32UK
H2YL5SgmSqz++Ies+2zeay/PCtKdVcWpbKh7/HufXApDqcQFywKnFU6L4GVvHwilV+cjLSG1yXk9
ptQ87DuTSzza50bEaN81m7cY/qgg+nepSq96n9735cREASvjzKJRm0EYCN6nSf2LnXTeULpp2GFX
lt29fUfap6VCtsR/OfVyiASXMLjU7GpFISSRTFAOBvFjibjsUHspiFC2V30Y+P0CSCtoWdTyNTd/
HcvfAeG2ZnSNtD5igAnCpiPkumRwxXGkC0jUQrfJ+4cCnMJyueQevqllpzxrCV7L44OB8U9pxI4p
rCI8TxFOE1YtWi5nzxABCKNu/StCiJft18NnZj8heTntMMZfiNhJLqrHxrXHf2sF2fDR7qUzCAzg
5lIzki0RRFwmF35DazWBdMKI/T1PFp75mbJKLn3mbBDU6HcTL6gZd9M/LOgyMZW8xnkI0J5sZtdM
Ckz73aIDqgkaenIzLdAuXdjpNFad/XpgQtmCRTG/si2BRsJ8HaCf0IfayJDmreVoktttT1hmIlQc
VKtw/WpLrEzLXfQ0TsTo2v+guvl4+atpE9gtmJ25Cj6tC32lbN8DFZ/9w9wkwkcInN5q28fOg9SO
HlV0ACOzDiNKJPCy7GPO9+zi+ywDI0odmBFs9fs5M5eZYICQQUZ6b1CXzgAvoj0pby3ZZdE3CWp+
LJHHquR5Bk/YsJ8ozsg9MYr6+Pw5J9zXgQVRPQhIAuFAORi2O+rozliQ4aJwX3u1MUWVSM/A/8nC
X7TomY0sxuo3NXyUyaJ0R0GvWKurultbOn9ThgTFtsIYG/rxs4zjPHJugzAAIsNWY5vUR3Ne/fnX
KoE1ytfGxnWhi/fKUpi2m30qC1F3D2y6oQWweR/xs4i6DQkTjxgWzPd4uPT+vjMA9sF5czesEIZr
h+2SQ5rbsDLSgxYJ+iN7FGgbQJ7SrmxK9BcQCA5DcaIA8jo3Y9QTpkjAJ7SW6P64+jgZ3cWTFqRN
jSvABbzhDbMgmGIYeoT3NvxeCxnGsbd4eM1L0/Paxjvg7rxVtZzwCJPn3YFu+LnYwqkUthEMF2s6
CXvUoNr0dKvlqtW9OHx7d8/d9+tcWNSsiIlzUoqkRIc6wdN40VXsT/4/L1PnKBY4k+CaWgARvDa9
nEvKqwRd9b1TwfZlxYeQKVV6t288xAMJgve5KhzQaOb/xyqKV4Rh9USNGkSflRa10u6o/CZ5yoIG
YLWzGPKzQ2daynoegqn+3/2rOca/RMbgxlQg/722Vcr1a/ObqZ6ujcj4VOikec3ufdY81ghLTYsr
5EpJAx+dxfcFf1r+30GubX6NLO4iaVniOzN5ar+TOVmfqIJg9Gl2RpmR0oXVKhoL6mtLJ2ZD6jzM
1Vglfmufie1vzn9Idrf/5ngr4sfpYWqy0gk2y190Oevon0vWrRkgA7LBrX00+RKkhKXY9vTLSEYg
6wQI1fEyC9f75LGFV/YJGysiLqz11BdhnfPE/p1Kmvlu0aKQRGeVzYT57aEBIH685gdNcfVIpGOc
ojxDWc/EgW9usTVxR91l2cYHuc174DzOHDa8hEvUNFFRBnFYl6DVroAnf2xl3/40Moi3J0wqTLOy
8laox4qSjRnEoenFJba1aIRlocNIsyYTuozI5et/itBLJhcs8Zp+xQYVWCmdMtwJXWrd/rHQr+/U
jcapQgKx4a1ie8lc0FvNI7d07xEFYRdEI18QvD92Th3X9YzWN3GOjWQDl4JP/RWkc2wQZMWRgE5g
hexUw4wAeY04ZHoI6xrp2H+JRfxrqBloW/Zg6lXBdp3UJzfZlAuVAY9fDsAh04lm9JApZAdYr/VC
G6OUt5uVoh8SUI1sYabLOdbfT/TRlTBNXNBoJsuVqWyFBYLpezZVWWKBYLmf8Rw4qQJpNz01TDvo
EDZeQmQyrbBeMuLabvpi1VvPT901/PSbVKbjBY5HgMYNOxzhXQdXJczcvcrPAfRJrqV3B7pw7mW6
6JhR/886E/qUjxPt1L+oUkQ+NHWeWXxPT/xjuUSyth3UoV8gFLqkWhUiCOPzhV3JN4mak654Z/ZD
ggOphAJBauunw1P8cp32QPmADh+GYhnUiYjghcmlEYUrYwYPcpBWE7xwEjNeYrTWgxuLO0Cn3FXW
DppXp+mwCrsamF8Iu+ww1OAuppmVccSd4Yzg8AsCPKy8kMRwvgKrZ1wH5JfQXZ9sUakPORJFkiCE
mH10AZoo8rgC6EUMgXPQhlQhqBq3lDpvxC0PZeyvWGYyHA2SnGdkZc6Erkq7S13mBWh0t9uXVa8L
dsAzLE0R7GVbJyQmlY4ENywqXxUcR3LoLwOXh/8HqscyB/gn5D0d3mlLAEEEF17aIx9iQ8baG7Y3
KZsT28+zAE/xYpKwFxBfiAvKR9soWhKwucF8TA9ulQsUDB+q2rcLEILVvLvAWLVvfWzpULBzmhQ9
K/3m0nUT3SmoWAx8ukuckRp2pl6pSz1NLoo8Gru55XxjinTLOdCQRMFhItX2g4MaNSLa3Ouy8yNE
Om/hwuz5enG8TREMZJpljwf+78LKOtw77M9RgKQ8D5r+O0IEA26dXTiXsI8DOcK3XtKtL7aTIrnh
JxUDAyWmqsWvYLeZ54hLuDQ4FjvsPZ5HkXz2c0DWdBIDb37k6SRQbav9o6PKx9PHE8Q6NewFKmur
NxkFNm2CMutME7fgXLTLhAOQrzfoqlnO4s/K6f7Kmw3N/AhRaEtVxdhgnGe4cAPuObGQEN7dV4rE
bc/GzdPzeiqmIPLzgvWq9101H7GCfqUct50r625idzMJcQRO1G+WgpC2AhAMmMJ3nC9QMXmKQUCX
4FqpnQLClbzXhpTmt7k0QbB6/V9Y57fxlDyB5Je7yjstIwL8wIpdnFKnzgeaa9U0g3Vhpz6wx6pq
1KgYDSD/z/vhk+KIJxjtfXaQhkebZfGMMrsn8HmSZ0RB75cuOr3idKwCxr2NrfTavlLn5dhXofgD
RnvYamdLCYezRC9OD1yOOhO1Bn89BU6sTKJjxsJaxA3A5arQKoZKEH/KVkECySETCZ7jUJrre87U
igJ0Scbi9cmrbmzCviRMdJSRIaxMSWJALL/0mTVxMlwEMVzXWQBFZW9KZncjOu2J43tsdfSqp8PP
LBj1ku5mCVxcgbu64HAj5gtkVlgTpZIJfjZ9kYq6i47AVjmA2UujJsJHbMmK70+7OCMTSQq+nJ8o
XuDvRDBInj1EYxT3HFUSbO44tRxC1Upp2wv2zcIlZqwFoHTx160G1sxwnvn71ItBBPWnmgb/iIWd
6lz3E4bio2YO5gXF/058lVbDZLSzAyJ8RYynTgQyVbWo0hylhm14BtGp1dom4OOAci79STlk0/id
0ZkyszTfSpGdH+TSS/6Shsia0Ei2QwDMLDbeyN/AIE36VqAivxf9pUTQei+LhPS+OrwBL71WNpD8
NzCwPFDaj3RxAwznP42piPwe8EceFsGNssnyzfn+xYHywTzuW9B28S9t41OzM7bXjuqvaEcBHwm1
EIHrN28V0Ew8YK95wXe81jhc/I+LNicpmLSe4b4Gz7dIr3Ipa4D0Nt1Vf5gyijhEbsR63CLJ14DE
WxeQigPXbSVoSz35HV45VxIuvIiA7DeWtq/pLMFftv1ep4TJ6Yr6tnJ4JcMohbl/JmnZhDffvjKr
JLUg7pgn3vGpT2Y3zJ1Ijz0mUXnobMHFte4lo2u+UeGd9MosoSrDRgc/r25wvPdci8X3jzhOFCVR
cUIn2mFc61UCw1S4w2Isd4o3ifQXOHHtmdvMMOQO3ITjqM6EDYYzvv1NbdXtka74TK6O9v7Q4thB
57/8bysrLEWwKJmjwL2KxGkPpOdDZjxAhDQTOOcbKYxJIU2LgUY0MQ19fxOtgWuEy92IC/sOCOhk
7HVV7B/hDimRBB/clVRw/zp6S9cmjAYlAkNfgGg/tqvDtDTJThjdNRJgj9CTa/jzIgeRT14MX+Qq
Wr4+cJos4lIC3ICve7dwjKsmJXr7qud4B6tRDtDnCOie2Wd5pXageCxBabQxtAUOjZKklBtRWZzn
TJVBcei/Se8YvzvjeOCrjIU2DfHdjpoGIY78tpv+AhpFIUftexRT1beIr8GB3Q+s8rbiu9EJ8mEn
17YpNL7h/c/ae5z9wtw7JcEiEHmdAukycYupg7vomFWLnrC2FF2zX11hEz2K0/0hnjlqCeCTdgWG
90NmF1UAmdQciVAYjaDzv5Ce52lM/EsuUQ3AH41EVZEF7tVFYvFT7Ueb0biFrih7LEdU0O2CRKTU
uWGBrRRQuxdIHxOQGHMJUUNocvR4u35tGyC8KLStodIUu0kA3v6G4FM5vONZo+FIjoFGbJyQL3mt
iEagJxoygSdvBe5MslOulcPzv1tB58uJoKXBPtcFh0VCrnWOUZXBVQyXTOrAGmk3dCST+UQuUIDb
TVVopMN6YLLsG6TCS4HpcZu8YFb8ieR2rxjlWfaCCOCRIfDjhmfCZDs3wXuR+vjzFAqwjoUtSK2v
R64cm4FzQ2+doADwsB3sQzDsoGDk+pBtk9vtQrK85b3hPEThwQpSw2Wm/+1GodJ4eYjelLlHhe6T
kmQ8tAM6en++qkOe/IElAZI0GTU/DEKas7VkT6Cpt0W4bZnPG71pfVZ9BK6Yi5uffEpkGK0DywW/
YpD/94Ex0JGmgfZAtujjqn64GjEaV7vXlrLlFOWEaVVVvux50iClktR9YXCR0gS555HXvLCjd89P
ZHhw1pJQk1fyutlDx3/yjhm8GwtUY+VoOZBJfSm1kbVXMWVhxq8u7nIaZv9DPZ2hy9I3IkACaY3w
hgw78YfyZnMukKRm9KIgYmEJl38f+uHVYltKWjlALxqsauBRlxhKNfA7bW7azNAc00fTUaIOLkEg
oLOlpGGLE64yVJRzqFJYti+5TmWTkZdY3lpp0hD+xxsGknWTqcjblAkYE8+Codkkb9fjnY5bNvCB
yaeOnPr8KBrIv7c6JurAHKDeuoRdlirWq8tKrvgZUvNrqHXEMF5W3M6apQJHxXPiOjKo01YbzzDK
SuAM7S1RNGbpi1lzewJVYV/TFSkWmilE/ilBkdBQFQyo4WCXKJkl1dvwSzHHD7/BlaPul4x6DGSx
YobBGkcO3C9ibp93htqAf84vg1h2B4HSpPgvTfJIyJj/bzwcpV/RMIzkC6e5LEk/FPb/aTwVkpsA
QReLEBWRQW5A+2OlP+BIvP2UKzkuAuEPKk6QGGEAd3lstK9OC7iE3cy4lZX4aJ3RtET0umWupcZA
lJQTLHh4QKevL0Bew3eNG8NWthJKPJYfLCVMH2tFpPYvfY1F2NKDa5DtYBF0//D5IMi1aAP9LGFt
6yki0nHu9+97tLhwdR6idmprSJqLaOFjbOYlkFWYUlk8fi1UAw+JyJtyhs7KHmIyTSKTASgxSRcf
Qi2P3touBNKK1OhNSjv6NnRYSom4l9d0RCiaSmu9cVh8PtyndufXJHFJ7CWWQbNfQ6ekk5mqjwum
XcXNbXrPA3KMu+rvek++TwkjYfkV+QnkL5735dgQu66AEz7DPdkd8T0+irq6ud5znze5h89IpqCr
73ge9+qTMIop4oFZhceB4BqwiA7YXeQw8aA1PwmxPC0zo5zHmSpK/w2PD40avu+48PI8LG9M4VTz
T21nHudMku8dLYzxqafUfefRFZrtz1/7HIm48SH+Oz7Vxzh92adLomK/GDJlsCvcb2LTdZANzewc
t68suUFsUdtrLrtav/o2wAJ//1zHWL/CyR1hQBG5rh/0WBJEP6dUnxQ2W9oFJ6+zvyyx+kktyCui
EiwJA+r3jzaUgyoAbWW877wrIW7dnkE4gJAkrcKiAS+EAo3ezAHWqlt8+QV3rLdsHEC7w3SfOcVW
ekRFb6m0efLs9v5HsElrQOYj4ofmHN8mQk/aZLsAxH80M317souXOTge+0ZRcl7FZEqNRg592JVT
kXDjQutxvj3pkZfMjPe29yMimb4tc7+sFQIf/5NEQVLBYV2A85ewYqb2Tstn/t4mNv2akOXmdXo7
nkvpXDqvJLk0WivJwzFSc2GsobAneRjVNJKdS+8+ipDwsmTQjOCIWITngkuGGqDB0Gru1gL1vJd8
+IBggwQSWLVOIKw4auWqsE2XfoZYfr2Lje17KVZXU7wF1+1jFD3bOAF2+uHDUBYEvvBbCBMt9aZz
MA308nBgwvFpghfDGDUaw/MERBW/HDHY39rAXq9qc9eUKlDfn0nKUlhNsw7974hwDvUkY8KpNami
SsWxtwIQxqpF1QJn9enGxSzoXRAl7xsS0WPaU29QKXtjR50Il9Yr10j83YuZd9tZVBSlTVVQuc10
f9VAixKvWsPDHapcKRLFwYmXOZk6VvWR6LZ9vPer0GWqIqsI0BxRecY/fU02duEs8ufVivMCE7Hc
NihDJOED5WEdwCWAinA6kCA+ku1//bf+vTVsO0jzzHBAqxmHNbVdMyXmZerz3lMhE15EkiDyiFkC
TEiCN38VnrHZFP76/MWB4EGp8MQlkeQyI6PM06lpBMbFFMyHBlA3jrtWXvdN9Gb3w1XcIQtWnqgy
SKp3uj6xv/4kEK4WdNggMbYSaL7GiFBghcT5aPD6/MHAnozBUbChuDONtJk/MXFce6WsT8hyjt+D
6sJEQhZ9zq1IIyH+UzCyVxd2wKmdJmX0ViNI9EezLQzZDVPIJPBipR0vPdTh/N4FwOtTK9I/iRK/
R80AgKigQo1dMxaG4lAtwFKdYzKKjL/WUvr1aDxAe0VM/TFdmMSzvswFJXuMiaD5pFPu4xVFVi3D
ZdVsS/aw/zSwJNj5Fnul6DYOJMJ8OT5Sxf8ITngQCgJCUvKEjyMFN4RB6PJRQXIj49jqAIDkzvCW
zNMvo/InSxaanT/sLxJWv+nk+aAjB3NGtr+2LgswQeQn9epU7oA0A9YAzf8jmICxOtaV8Syt1Z6x
W77YWh+21EU5BIvhm3gre29VGbGA8bZsXuAYiuWL9j1ZTh71c0zgccIgnfsvOmnNPRBRdEoUfzAw
Ew0D6e8BemgaQBifOJDROLdYvsdTcIWgOy7cJUbuPDH0EVsWPCVE0qZXezhKWhmjbzg0wEwnu4I+
ghQXYuvSNcBRvpqPW4AUcsqr5hvqoNqDkCeGDEWn55AOaLN+HEjxb78ifMUpQTzqkwhMvhP3tmNr
Olx0Qtu8HNMqP1uFkmt4l0+XT08DciuTgsON+pPL4gmi5VeJcxdUKfNejGwc8X5OC7fMTgvF41Nf
EG8yT6AEO6gV+T333dQiZpSbgMAyYUfMnY9A3Dhjd6zgiNpyq2/7uf2xNll4fj1APzSYiR3CRblb
3nhSkT90VAafbUPTaD9T1Yckd2+UXPTe/quRCl6npEJ52gwZOu3LW3Q3a12jWDA035alPvhKhcC1
zn/wIKc1NeMRkFRzRMeK43c8P+vAkCZid6SiWf8+jPhtjfJwI9IlaFN+U4XwvrHcmMTqVqJGslLx
IoNOycl3jYoJIPDEvVcgoCSZFMvCOj7NcBsSGh8lEhk1TNV0cWw4QC+8PfsSZkVFUGbxWKPrzYib
Kv8jA7WOUlncaokL6OhIE9CWP6RzlhzPlklX1TxnEwO3wUd2O7vFjFsOiBtU/KrLjfs7Q5xcTkx0
RtsGw10uXY2k579h3sIF/4y7chj8LqxW1+07jYpbGK/mc5tAE4HnD6zpi7yKjAeIiaUybaCK9J9N
kM8G41ZrfQH4rlF6VxXwZYDe3V0J7dkskP389QSapuMrFNEb+egREzjXseH6+ccdpoxa3hR2oLfO
Zzqbp3HG3M1+DCRFs4nlYxv+Th29qu95HGYtc9tcu101Satt1d1BvnhAxj9CToZEuUlfIVqtImuO
M3EYCRS98U6ciVs6f3JNDEEH4dF5R7l34KUhCCV7Bk8PwaqfQaUKpdZugUkWbI9s9b3kWr9q4hiS
n8sRBWTM0tef3RDoP6FS9iUI4FZ4iKSBiNeLzExmGZwB04OqA39t71Zkv2WxzUNQ/4ltvi0b8yI0
JbVVWWBmTXBm5ep511VW/wwv56zrXRVBWgRY8Ea5FkqsfaE1zfMHAKLXMikXjL954p5H2WKieusb
6LpuXqCwgtXxLQXhsPj/ZFXS1HTv3WRSDhSVtcGon2lx61ZBBKsPb9KBZBV+KI1JvwlaG1zwG/5p
kRJ/mGEJ0p9a7EOaScBpiBXNKtGokNi+h3gqqw7z3uU/PBvau3NVmatEFuQooR1wzZjkTEl3/83a
tlpq6HTvi/NftXGajZxtoUVdoEwwJ7KIQ4pR89TEGyDkbQ5lx1ATqfzgakJuD7JOw8h5+rGs4UPs
9ScI0NewTsnitKmOvLssbE1g4kBvG/1Ja9xPWzSqhKEXY5pnCUJNiUDDSFYAWZ5Ka272Nkv1zOLq
zj6ZjRRs4JKupWHawqIaNpMc5NSOyLSV7g7v0sE7JThSvgQ2SlRZIfg5Fyyn0vGes2WflTUJUPVA
DJ4Kb00sFo4RNEgzYA+Z1TQeXtbN2HMCowb3J3rDlSPt9o8ljr+7vbQvBroAAllkzm8+Z0+ToYeJ
IK+0qEIl0jhdnnFHBe6aAza3FsXHKnBYLbbPowa0QGlJpDmXlCWq/fHHSDKvy+KLHscKFU5bt9al
blDna6u+eh7HgdFeaVfOspbzK1nmIYfZlB+Yil4g55ncs+szzT7kzx6MtB6dyOwDqsDILiKoenPn
aQSfFaSEjLjvaq3MRgIgg+ujwRMTD1l+LT34UxX7PHwJIy/t52SWbgPaazmoNgmeAzItwIrvBIry
C5zqR1elpWx9pcYqPs4vSsifYA2J+zcw6yWDjRzqNl7YFnr90ZQTCMlmWM4CcL6PAI+Z+3wATnIE
OVhoL9N8aF4XyKfqeETJY1YKhzJV3VSFZ7PrJrhy6uZaNSAyGdb5yGnyJBqzF8IjxV6Bj370iQmy
5YKtexnSEvbKZ2gXxG7kJV93phDUHf9stRNZllV8iLeBYUBZoszJnRDZ1gotKiNh2BPzBgtbGP+0
A4mDlJPIePovjNlosQHmLEL1rk1y1JbvyNk2pqSToUJPq8JWddhNPgoLm3/S7Yb9RZZjjqfJ3uxg
vHooYqyYaVoOzKvV0AwEajoD0q5Z+nL1MbH3Of/lzJwirqv8AdBLpi2b2FatG5xaTKTLe5o9vULr
NxVwYTrOBnrwP+CRKqFUwuPjStjA527GPybzy0l4RwUx0++ou9IGHxAF43Spv7a4Gdu2p5yuZpmZ
n13F2IYfTltZrqQUwHC9wQU480l00yJsBs/V01MfCXNlFavgv3RgGd5rULDaTGVuIMiV0NHYhAN4
bDZK9fOIoh3ys4AMHSteT0a74QjVXWvDPhovUx1xueudoo2qWOZESvkhHNNWtYqXpB54anf6upPw
e6YCuGqF3cTdnnzCaPoOjCX/DlK6ZZE2ANdzN6OjEOGze3ochHp2fHsHelR6I/i36SIrC9Qhu39k
6g2NZt80oUYC4w7Gh6tjV4Q7N0khxMk/BIgWaznGq/1CLZrw0v6NIN1ZAib1rl94Hj9N8g23Wqvc
f1yMkYrclC5p9dVxj1w4prQcbtK70firi9MA4/bZcnEUnKcDcdgrjX3OvmpL4IJzbKtAnS5nzp2U
dDlDzE8269bDsDXB8MuSxjH13P6MLbWVVgpkU4Tb4vb/J14+3J7WPBtH1Ul5JCCI80i3cZ7DyM0/
LvPMfWBCWpJ083WmstTWdTt8llNAcx5NCf0aShzdqR6VmqmGGrWIumx4/6jtJ4tlLgK3J1amQ/RZ
kVmsQGEhxzdAI1smBfJUHIyDDraswN5iTzxiC8tr7cD3C2BUtoktG7xtJkpOfei63cd9O97IbBqr
PdwDw7qHf37sKOIw0cdtuiz7BZJGIouC+D0DCgaq2rBVyIOA9iaQAKaLWHOUNzSzUoagWUohfApA
FOtmc0/FclytqqYDQwevGKzBH18F/p+/BdaUbVS6He8iP7CYKhqOLcV9cB1mSqsTt+te5JhuswII
CKjxfHnHTthExJA6DOWihOT61P6pIeaQWtjIn1r4XqEk6CaswPd7rhWY4IclOLDayAUZxWgga5rk
iEepWFgjk+La/f1znpupKfHBIVccfXEWSu8LddU1CZMh9bVi8crMkgSzC4ky2ATqNibW0WfBUdIC
FJ63hxyJeYv8t0fzs7M+z5VHEQBcISjHvmhgeSQZaaoTwa/+400lgSVn4tiBOn4w/5yQHuaAfKGX
/fSNyt4CjN4T/mVhL7G21j8tk0Yko8OY6TFMx1BTu6SD9PPsnPb2tIwx6ZsC7FOoFmZ6NvFqNKhS
gZO2hBYXriHYIJVscQpN4Jbv7T5Qv0ObfUc4Y594zun9eFs2RN+UpR0np8xUpcmP2vPZU4A5Mof6
BlziqmJLMF+8hV2Qg/V6tnCmLSy29w6jnwEez7ot4M+DXTPHBzV9DdJcnxY3bmm+POjl/RV52BTF
V8wZJRObPlLNftKFj4aMUOEEQEQB+rvvenyvHXBdRqBe103mBIX35nEc6H91xxFvsd40xXo3zOlX
T48IWyik+HNO0hujxvRaV0PbN2rojD2Rlx/3LXaP9mhfscnCntrs2rmjq4xJgXhb4tVaQhSqj+fW
jHwXWKdpw2HJcmXOfYcZemPtdoryK9V4xGsQyk7aMrjhPrpG8jAZaahPWzC/MLNlcvt3PJbspyNM
3Zg3BRuYvWp9DFO79yj3sGY3eAb7iW0Mxr0c6ZRR0sEO8wSnRCrdcCbygcAKaXn7hJOwi9SPEZ22
GhNXZcs+UycNioX/5E1gg8uLqsZ1eluLZge+PbPTCCEPqtFaJBUB3FJ2VGZErh4L3s8KWEKRgvvL
6jGeP2k2WsOoP7uxa2NJymX3KiPpL6UvRGZOGtzGOInCyN7yvEXeY0hyWtajQ7HE3Wswb+Q2FL0P
vEHIoVV3TOprBlAQt/a9IPHH0tbo+6Wt+xyLLGhWvTwmvYESYEJVnk++GavjOmrsVd+MuJJPBfwi
BYmwQixzPIHjUSkEoskmSesh0psj9Rpc8xBBVMcOpwhnN5kEzS0dpy+X7YjJl/+I11Y0DDxQt/7R
6cmHxlYij1nB/2KKOXCepVpCk8qZeQ8WDn1q8Ol109agA/A1P4Z+laiKWx0CH53DT1l4O7UQDSXy
t2W5yPTYWsdpMVLLSP707h8+kZvvY7PI+LqV/l9LvtRUzlWzwtZOJykTYzmFiHtNmyCU2MSoZqhw
+vIRgqmRFozQPPHABQvKmyi6W5XMtGYNs87LFM/KB5M9sQ7YEHuUFINToPQmqMJsAVHWe+MvwTki
jtSW5z3aOnYHacZ+uV/6oTRzE52R55NbJwWGsP/SvdKLtfffh8ljmSRF02Amn5kOfM1cYkGIh56u
xdqRoyDNaCr7pI67pElfs+l2GSYZzPhfaVB3RMrjv7oqS3/OsxEGaqHAW58B9DmBYccurjexK7hn
UPLzM5CH5C8QkheVD89z6fg1+c1dNhLa2rh3421X1JGMBwapD1e8iehwY/4YZuCy/UOqiCFbaIKS
ApxPCaJUNEkJY7NhaMGVEn/JVDqxyfXrIyOlgEAXQ6XiqxCbgE8AlR4M+qUMRXHGm6lrb4YXtsft
QvxpUzpczNbtRK30l+mUIALRIWEVbripo8LnhkLTPzu2nrur41OP/8LbsRFqh+BRJxcTh9AxVma/
Eu731sJBETqfQN2a2l/feFbjWkposR7KraQsS5oO0TGrWi02D2oruaN1PKb267fr8ZNhm5DvYRav
Eg1NcUzCRISKCsDunlHFxK3yzqFLauazPd3Vr8fpW/97xYHSb5PJRACmXx1EkytWfFL2JdHKwKMj
o46WqUpTqXiU4gqePyxNKRZoOI0CB/ygHj2OuYgLapAuZXc+ze/vjeh2WdVU0cdU2Prigl2umzYz
siyV6S6SxGLqIQerSJ0xhKOr8HTJrXX9InJT07GykU+8oe7zCPUWk8X/5YKaAgSdYM0SWy6wAoVe
Q8qvn+aF1WQ91NLfArzqgcds7d8S1FMOURIAiYCbSQEC/NuiQD+VNTX7sO0HWE6jmUn6+SII7/Ki
JRngZ8K05USULUjsR08fhfNslortNS40by8ufMTbGMdw2L7Xamd+g1Y4foQncIvrdK7B3JzNsPLQ
kK6WbIr6eA065SjA2gvvdKQnZrlamnqRTZuuTRMHjdO+ua651dQ9t4KgSERdvmkuZGcATukJPnqn
0TSdHgNY2AYOdAzbMhGzX6JUUamZHul67CiGfnsA+XXHU9DhVAbM9SmRb37PMg1bSXURkgnhPMHS
8mnEwQQSazzUtuQpIX39nO5FrGsB70RhOZ5lXRUiyuo4gOYbvYQxz5/FvbWj3lmNSo3ngH+E17pO
GWP5xnDIF0W/bGreevyzGqx01SuSvUdBwpsObZ35kWBlyLFhwcguUHigh8bEoC/c8ZNr6VhmyqYT
dnGrujoJqbkEdjKmmBd8ztnOcd/6Tr3Tq6imPb4TpNGCt8be/D/a82Nd9zkkR2plS3DVsYp18eYd
V1KiELbkHj+9PL6/8deiZ/+BpsD3PrX8Foa+BgyNko+W28JKDatdkBG5IneAo4VkkPOMdv8/z/zo
a5Bv+VAVZ0BRRTKw1hn7AcPCH7vGD3lpzg7DhPzlcGUf9+gG1eOwmNeLJ3IpvguOpsuZjpVk84To
W+7TuBdTHAH+b4HK7dP4DlxoPLNQA1X0QfOOvsdEKs8e4ZEV8oS6UveFgk/GtbSzAqDD2rdyj3Ut
jHSIbYOH7kyEzQB3zDe9mdLGWXebg+o0iophkHCL6C7OFiTVwXpkooiDBUpgu9/U68QVQ9GLQo6H
JMLh64C1+miIlcWFV0YTYqP0n1QnbmBzVgwmWaF3fZZNgQesdx1NVDfWTwo7psO6JX85ZkrDZbLD
j0bq3ozvuGtmlxXxrJPTEsnTbSruZaGbp7JF6OImGJSEoY0c4m7QnP/UKy3d9YkpCW75MkSY67V1
ti3L9C+aPxTRxRPj6asyH5Iq5xIkadTMNGrFITnm8Lt58xPpwajwqitFYAVBjzuKytLyKIC0+nKl
w1zQSgVNQI/JspwbYIpSbdVObWq6SEGskcljonLtsyufxIBl0GFrWM/NrTtlxFLoXpDedCRPJdLr
wrCGxR4QMjsoT/pb2XOTPvz7btrZWGd11Qo6NHGN4TeCgiU/sgAaowPZjtSXdGtnhPssXvA5ElXv
udjKgtQdwXITSkD64iAOqu0Ppvbax/1roNmWKcE3kAlDbAowJvxb2B3ZFOdPEubdSTGIROKHl43x
cTXDChpm7Yp0z1+JooVT42fXH880XPvlT4YEZnUPQHaAOY7BnBQVRxoso6ZqKK1i6X4WrAOwGGvG
3yISHFYTj5H1rv3XAZEr/+VzpUcKQuAnMOfXF0Z3uhN7F4t8S9rNn6lwplPSWLZE+ZNhX/1vPS+Y
8+XLt/NZikEdjksbE78guMbU5uMaKagW14WRKvy2oiEFTzf9ED1YVLDwGra5SFHNZHmxU3W0vDlV
4FzSQpVTJlFj7veZ3IR7FZHOCERklQyl6pUR1x4l0j/Pq+ooLy002divtYH3PnBxW5evoXNHDpTe
KdjS7BVF0QDYlxeD4D9RphrssD2NYeFk2i6PxJRcetOv76aCuBhTwd7iPPaf4FjtuCbS4zptLkUZ
vVU2yMi6DQhB7o8LYo02Sx+l7iI+cnddaIJ0iw4F/d9URNxOKvmBdK7afpa1TF+jOCNvngIRVdVf
XxbtHvB+YFTmq+XFRc5E8C0XHKzabNTHZp7im5sIj+0XNrsbp4yf0WhzE8DvKRIr6LQenj4u+YGA
oOLv4xHpvH+LXMKBdfitlAjv/iTCclOIEkOfleO3rCmcyDdBDlSjo1vU1nYbSEGXBQ/L75wpv6vQ
N12NFXKtVQ3majZPt/DK5e1a1gB80GyDJk2xDL9UvISDHFHJa7GpyeGYINgqV6CKLFX/5MQaOGee
PwtV+mwbLKlCYSFI4sVIooSyat7phfMfzC4Ulk8moy3KLbcwxGTdUhCvbMK/CtwxA9dYfE2EkYgT
8OA8YgeBmupPX2dCu+lWvCokZakWOfaWH2R9NxT2j8MjkzR3TumfxF9qti6gy7e8f3ofddSLqMni
Y+l++sDftukTS6M1fsaGggG5Viy8HMDB7wUxvbFfvIEof06krActvCsDeSwGbadG/sYDEFZngjRe
Rx3nLor3NJ+f1CGp7th2354k2D+ZxhPPpy7hE5wjfwwgAH6fmaS19Mp4kLbCksvdfmkpeecP7r1a
bwxCg4iP02NRacUJAFE/rUn6ClC7+NaUf+kaUiob5tEp4pFcRVSR3/KUGvHQ/wNNyKA5PHUKDzXf
h48bCUVyewAhJcboB7hashWTiybgICWBRDq4+P3O/yLZvT0nHUD0qtYbSVyG4dEAfwMdJ9LFDdJl
OYaeY6vEm1/K7gme8QQSZO/4BkGmqQUpQjfweuOhf+bPzwQLdLz3ybuHWkbstjZSSwPg23JWGsYT
j4ehpXU4vf+4hk0OFuJjwWgXQXI5vZNoNfhgZOMaipVmw0j/N8oVJzkOpAEloRR7JociMSLqXHM0
L3EsyjEoAT74PQs2OJsYP4kRuVBT5kSxYZzXmkYQFF2e7+m3HTb97+4ROKOYPCorpqRDQJOzPQQZ
y/1/rheUKX+EMaIekwt8iOjXyADQlnpj6KBAyGnW1zvq3j6XPZiMmlrkT7hMNEKTjlLinTNt+OW1
whb3ltrp6bd4mDtoM59RknXSgcWRvDO/EXPCTbfh4qXI4GuLZg/oleSzvPwf7gKZVlAjZIMfZP8L
HK6K87epK1k9eWqQHOmKx/u0Ec+lDuxs0p6b8EkTBnigkwHrYqJHVgznBy6m68PQs1O7T88RTbdF
85QR2W1h8jU+kRIKkdw+DmfKY75CmWGTWTkH38CVjsoqgDkiMoxUe9/3iuORJMv3Kvwa6VoceLtd
IRxbmUHwsyHxbCaoRyUo/1ECjZa29qMm3FHwRcuaIHkmiSQhvF7xMVn14IWIve8Q+0qX4X1z0IAk
K+Tbh9N3WmSjxq+/SjQdOanlbw8esuLopCGfWWCuqch2PcNg1+BwYwr5r7ICvLxBDpVSIpalvpUS
hbg7ioyaLTB1xK2vAsehbpyVnbq+73oy6sWwWCAzNM+S/4V+512QW93H8icnnZKLN0aKD9aG2EZL
QjZpHD80YADLJ2u7yExpuCq7iiX77lL37eMNWwZbTpEZ4famHooNhOAu1WmkRwAx+qRbQfzywUkE
hOaKJqmC4Zxmdr5i7BmjtAs8eKEv2RUiSIsyt3vrgBTow5XiR8w74MmoF/rnv/dozUgA5BXebGfw
kLvNnpx3CBkI2bLgAhQKcV5CbB3OEpPF69sLfpVbxxPuWH32X9bcd+WVLpPVGQVn+wEBh+bEHiY/
bOy51OgznyYKp1kSta1Sf8E5qZuGlpsm+oc2lv7FvYkb6CgwaJziddksmSmt4+5T4I/9qnxIvg49
Wyt7aerjfD1IKXVzVue9BaqeQVrkhjonKkLTEWoNEeKWJii/XdpARM0T4f2GEtvfVN00IIKI1HXw
BrOB9ushDJ765LCu6uKkDLn3xhGceE7l0OhqZJks6+pEEKh54YNXDtqgP2XIvg/SRS8tnKRRj5M9
KmByqVco3D1hV9dVzuVdvqRVqbHJLXKr82KvD4OWFx9YDmDuDIGjB9Eum55GRKhoU8eyYR7RF8QA
b5jJOWjj4gYwPrr25IEnXkRtd4VtzSpxIiLJv772sKfqZpiCnLkxD2ucGXx0xiSTPISz2wSPPifI
dxopopMfqTyc3dJBP0V07UiQMyYD2q1K9LCkFC1zsE3p/iNDwQWf8Y4zveB3s0TjTT8UXz9wRDW5
kgU+7vb9la5in/ssCS/bRRRaHMWIFqNz6gaHJBE4I5rJJbvhxVRkVzUrUG2ktRH2ZHWhrdJXPP8g
Bv/9WXiDtKtnFCBI562j90AUjMhpSymX9He1I5SU9AT9/t4sbxwWCOSAOZcWwFDbET2mhbMmk2ju
5+/4khdn4sL9511I1f5awU2XoGIuO+RD0YVlXfsw41NjWwy1PFbPpd6cLoIu/TbmhcY4pARZPDP9
ZGXPqlxSV28/QbVgnTm5S3moNUlpQ6JRfDMpFzBCBg6EKRL7YdEO730N9CwQwIIQjF2blNq5U6Vh
znjrhmke6pvC5p2qwkm8wFUpOMYYbFEo2e9TZMPJGkHTCotjz91hzhlTYhv9eyk4dtvKvnpUzcMc
5wh1MjhDJME7WYgBthasoyaTju2d5pqJa128EwrCT46yM0H1ccd+Q5WFWmuBNB95Q+UdbkR7KaJP
ChblWDcOC0sGKnHxer82wPWlbQEXimdDP7NcOudKEOG+08RjCXHN+vCPYZN2kvjg+6aTE7NCnnaN
VeN734b2Joz4c670RQrccWUapZ6wFF4ldlhfCF1NPShEyrw4Hj9Aw98iP6WxwoHDZlSuvNdsklQs
Li2aEPx164DnmoJlevzR8dpnG0kHd7Y5BmkFSktCbjvM70GELuohrDUTl05g0m6I0ROSRWcqpglc
KlYizhY7i7g9q1Asal4IYLLj4lz0oKnkt00W9bYcxKaHXE83Zr//GDR09rFc1/CBSQ6RVk/nh+Fw
i4x4t4mTwnItBsbMJCmcuvw1sCshnhtQ5D9Yw2sQSsf81fBPKHUT0dFVLREKrITRthR6fmrE8yeV
qIBf7z5OrR/qVquabOqSOQoYTpQsmp7YM3OzEJQuf3fNG148a4wmZeB6mFQWF4fllmL35ffT9QcM
Np73fgPt217tEUt+m4WWX7r91YpKypGReqOdqMzsuTsG6wSjcyfiOs9ILGgNwS9KdPWWb7FUu2ul
RVKyjtm4o5A00kBUZ+fXhyNhp1KSakIWaqJ0rWsGVxk80g2dbkuMJ4iDu5bu3oXw+YEXdJmYKc3+
Bc85mu2CPASZ5vrb7b6kLCh+ERQBy8TzEb2w0ruui1LHHf6taEBAleAHxGuWrBYHa37LAt1Vr9QM
zIA3IQwuoUpk5GwDLpSLI3oaMbZLWgN72bg4wNlum61Sugr1MO4CNklPmVum+q0Um5VOWlnjX1ya
6azYhWHtVHaQqGLsClxMDVFxPXNw5p1GkXLr6eNSl59+N0PCuuWnmNxRoMy8+78DDh7KrhVaExNm
WCxwRUPy/8wUOghrKJlgljWZvFaQYTcxuAaUz94jxVOxJnMj3W5gRzIYbs5PZprAeGDA+4nMln35
yaTQeLMiwU/sTi+BScV5+n8xmYhlZ42eRazSLAYGF0FMh/giveEfIy289pM9E6vpojRqIwx8MFy6
uT+Xxn88wYYqZi9op+pqaXlmIiFPuW4+C2YGT+0oIkHCuUdUN+/FwRPxfxuNObW1D7j6YBfQ28wp
k+Xdiy3R/CA4yXmA3CRzRnM82ZDntX6oMo4VQTKyfPvjsP72KsQtmQ0fPudxXjZS8KS+OKfKYqWD
uDNEO8zSJ25M5PiBtvLpvCMk4mAZ0L4aDwtY0HyI32c+//YbyhVn7bVFOUucAsWew1ICJ9mPKBKe
ypO87hM9bHbV6g8KuPRU8jaGYLmBDEIQoC8/Ooj0e4FKDIbcxupwKUpnyswh0JOXLggJ+HQXbxCc
dOwxGIg2VSIYF+t//hNtphvPSxgHnHy2uSap//hEMNT/HY+fnE541HMqc/bT9V+KcT6AcWFj7Qc3
XR1fC0uxCDLg+qWYwOdoBa1GH+xzKupVXrPahI4ALlx3J5P7MqDHHlYMEdo5Mxrqb+1rrITLFcxd
8EI2n43TTdPN5V4vY/Qo7JIBFZ5JEnDD+a5QGGbTQp1GqHJcxv+8g43D2OKrSUfmlENDYWV6LI9C
WHQiTmbgeQaqedzKaZxKj0GASgzaPPEJhIUu31kNZGNicuxti5L3IR8yxHWr+sSo3L1B2GkHXydv
DLJLENUyS8diDh3VAbjoOAwu7F2Oc6WL+7Jbsx1BzRKgH322EMqoL4pEd61Z2XW4hBjOUqKAHKk3
EoI3/KymlN9tHKhRxmCiPGyRoh4UzIoBQDiafv5VA7cfrFzMRkirmANLocvVDWlv+v2LjsftyKK/
JKdK9A5dPRO7MKcI8kniq7Crmbmx+XlejnNyLH3i8DqCfFEHJULAVwazIhnxNB3WxtGI1cwJpG85
mEt5UJvcDWh1BxTQeA/JAbQ8HS0XA7Nrv/fOFnRe7SynSfksQbRvyzGE0/y8lC8FC61h081NmHJu
XilBtHr7yfgUrt5Q6xBqTsqsH2b55EPNxL+1SPUik6n5r6lGoLUPT9L5HmaA75qiphH8GLRPOYA2
ke2mRaO8s6agFkLh8VhZNcw0ou639UAOcw7sdPN5Zz+SfnPj0Gn56RBNvJp91UXuqqOZHYwS2+iw
ontHiyF4ZJao55hkE6u5xJFLPeUflNEJdCDHiVG5wzgYTsbnaHjW5wO3AWfXbsO3PCB8gkrOXEyM
JMz0wpYflfNh/RxMhJzTgtVOQwgkSZ9hkF/ByXrfwqDijqZhctA5OBFU/cDi/f647zM6C2Yw9QHe
W0k95lOU+LTxm1684v5n+WcQLOQDcX4lKcHV77scWJBfkWSmWuhn7m33l94fsnQA5YDrMGZlvsP1
htYr0+geUNljf9HZFeiZhCgeoJ9nHhcT9sfucVU++uzUWbuD93ts8YC2GxlH0dWdyzVKJYwg/3Pa
uJj9NZq1bRw4JuRMsDdX76jJdolkzq/jDZnjuJ4Df+VD/W28JRvpweVNU9geORwUjWrKSNBLWY0b
CqVj5kReeFvJA/ZgmBwyuQnob9n2ubhiTBGELJ9+eyKvB0X2ejFkjZqzXfas4KV1JBLoYGQK0pm4
TFRlrulYKPn6686fgWkzDaWlqjlJ3KeWQ1yFVlKn1QQfLuxo66/ftCsC7l+ZmmChMkGcpFKIowoz
OrmsGYbXda8U60a0ky4yev4LhxVzaRWtliiFkkbs6go+e0p5eKKwulN/H7CAFf84MBulAszBUV0v
7mSQTMC/etj4HuLHNBGE+D0N2JnHS5/atlx29hrgbQdMOmVCX0e3UFPFck227Oeca5wCbTiFbjXx
cIukQKt6stPiT3QC4j5zZHlII6hB75+qWGqYN5oRJ6ErwCjg6tudwNZnvls2i855/OEr5APJofvJ
0UZrqdkNQ04iTAJK5mMn+k6bFisZ/SK/D1h9xFr7P4xqmhnO1SRgsncuc3eeED9bGHHBjjNzTwnH
OASN7RbIxWZNlodJwW1KtWRFGPHJZ80Cvyt10zucOW60gxGTiRzhsnnHfYzGMLpxghj3dPGeimbt
zibSUGrnQinuOQm0rRKwC2q6VntCSFh+JM+Mdnwz8hjeB2MT973fpHM7k7i4zRb1P25WRTlUGLPn
I0RiJZJgGKQSFGKPk+swcS+B/8IWqAcR4ZLUsE2Ubuu8YWdiAeN9nR/vKbvQTTs8xZ2e/0CVQvie
bMKgQLYqiJ3YDIpzHgzBXgwpBvQvV/5Gob46E2e1YwK6V2yNbBDBau/17ibbOxvoV3xHQjn84KK3
mlYiZMf3hABpoCAYWQSaPW5HKS727Z21m2biMzGTA0QhwjRN6bMPD2g/KoGlCXets7GBUI3IdFcr
DSwEDQVA0isZEnZ+9WatpCuHErtPDFfAp7GaW0xVXVkmlsoj2vu3EVIZuufRtem9/2fGsLH7E8zk
cLjhdFpy0UF0ttvr3aUqmlSn862J2D09WxfGK5AUu9qP6wxW+gegnGldmzjP63be2bGngvhV+OL0
D8gIyoU9vF0Iqd540cUP7EA9uVle7ukM+Tiy6qjskVmrjzdwJE+/3AcVHhWqeZWMlxDuJstbamy6
GIEBOgfW1OuYC5Paof8rOzMfkQXtfiaqO8wB6ruQcsblZWeJstmhw3UCAyeo7NhLc+YDDEZOMEDP
ErTLSa9s1meCjfbzvkiYxB8lAMlhIIR7LC+3lChmemaNfloU4GJrmprTOdmAWjIQ0WwxdeF2qB5N
aMIOnxyKg3/thWbjftItoyBq1S2DdkMJXph14XFRg9/AWp5JeXMJjRx/m3nVBEmdl1X8xT3qJo72
o8ZEO6g1moo/lPvkaMDsoowxN0Yp1933+WS4NvzSHPVwaHJ1QMvdaDAL1u25rvHJ1ZDhMF4wzPDd
/EhX92YF9ZNo/MekLzqNsUyyWEIiurPOuT4zAUSew4u+FBIGQ8+jdwMLhjPxWBTVIi4cPb+vwmyu
LLhQyCCKiESvezG7NynMKqJzjaiNCrQoPC17+V5Kce/crVar/DBll54RdTzJDIvCJDOgUR9iTNZ5
CkxH+SVBLWVwZF0gSGf9fRSjJJ/xetIjfb5gOZViJDWT3Owbd5x3PNONrNPRFgpojbojWZanKBs+
2O+iM3+3B4bb3Lui22uxp8u5lX5AthtE4OfrwuROUr3vwCaJaQM6w4S4yzx9vXY+OZbaxDPkCMB2
d/AOnizdq152KpyHrV8BuXJPa+swNy/i+uz85WDg/GMGr6ITsN6BsB5D8nWZ+a3GjehqLPIq3df6
rF45KGSXk9gq4kEBI4JMj8yf6qi93ROqxZgMwFL2W4njALug91QgZC8pLWjsxnPolA7CgUFFZaSX
J2o9AUebqxv1qdP0sto7WLSRtoLxup5Nnmeer/WW8R2bgPY7z295VYcwqNxTcyujgUoY02FGs+5G
YNCT6uc9DG+6i7/d17K6QlH6c9l2d7yNUZ545+0rpA1wKTSHT/zuMxRjBTyRE8okenbx2NAeX82m
LTaYQCinBXySs3f2mo2dFoPJXASvKjXEWY9rntvYxdCR8uSsaBKVGJvS6gV0LZ0o6hYK4VjSiXjj
Iqp9jRWLF+sF7yOrn4lYU3In4EFhS5Sfkh3psin5dSXYMZZKzW8SS9/BvD2aFgwIS/F9vbJYWIZi
QQ2bngpltvh8SugkNLPEwAmj72ip8GsYkd2kbkGgzAxhiQ3cVTM8IFyj5a8KA4ZNYkqFMFiwBBI4
vvMOYnBxzGvCw8cqdRDEtt4YD3R88qPJQHd2pgKS/W1e4mvh2yHuPciErcJtlkCW7tS/zsiZViK0
PjGFfnhaXD/20GPJjYGs8n3gaMfihb5RX4B8bpHL5AXUGVLFI5yJ3wipK5r/w8COOeoxnYg0ysGJ
locDwT1zUhnDqxVrgoaqLpE3/+iPkFpEgkXyF+4cgTSeEk5yfdjOj3uy2D4IsVrGkvtyglIhC0Ay
SDuTZCIYBMupYhDsoRL+AJ3iC65VEU7Z0+Jzl/ahiy7FTY2r5bvgkpASLvtjAm6l111YCiYCg2pL
4BSGd0CVQFh5JlT20rp5TUX1kZBcMKoXkCeVfGVXiudjQHTrDuPymoHpWAXxAoGrtJ6DCBuv7Yjw
7VkBvr3yDw7TzruRHXVm0vXUhTTxTmohiMbKptAjAblbdL7QuHY2IuiGL2TkekF6X5Bqm9gT0QKR
I+z1mZAl1pbV7DPY64itj2lAJntbXGhe9c1ecYEmOJiCPW3Xh05IAC2XIjmzTrIGFZB/bs8rZIPQ
qIESHRMO6mqlL5fTPOX1ImuUjo4o9aX0qxYoLhYDXlWcRNhhYeSLXlfqqgazrx7Qq2tcOf2xgZp6
wqGrb04/FYPxIHtYlTDihxWl9GzfIIucWuCyM/IdFLRtRq4uL/kVLXIn8dKTl1Myt7E3xxsvnA0Y
a2f2AAaPSskxnOcInF98B92fwKQl5J64oeMj1B+KTn3TkHighzl9WomuMUVXalQv2v6Hvi7u7Jsc
impv+l/saDmVojgh0jlLOHN6Q25JTXxpP8e8+1mguNjhW1gN4y6nH5Irn85urr2pR5F+WCvblZfy
D0yZkvQCsQBKVlvvLI9d+FiM3rP7cSkYc0sc2LpVkgcXYrSKXAnsVBFkcS0T/P383fmtGln2VoIG
KnBfzmWSXRSWAMqjvyqVXaF6jMyvhK0bv/hEmROCljtwU97DBEa0tFXKaKaUW3C3nidfZYurtcV/
ZiO59QKl3nDL2DcxcHbMKi0kBn8TQ8gPXmsI96Dk5GW5SgjOK7AGhlhtbwRZEwazumCAW5tM6dU8
aE6qpBI31OBwVVq7sDSy0hn7ngQALxW5gWA7ZtUDf2vejRpv613KSrtkniGQfcOrA7VqunkjSkEX
pA7mQz1aplUI0LBmAmtV85I1FIq2vt/Y25mfNP50e83DZhsbLqvwHmqi3mA+Tgw/0nTH+g9M07ee
CsTUiivbl29rY7VRFdF3Oc+33gXTyaP706Wth2PfNNMVyEgMH+s5DmWNBu6RD3FuNMCPiO+Fz4Px
zsoEqkoF70Zss6BmxZ9s+5mCgGkZv5Ly3OztJD0ZZuBuRqd2+GQg7pyf5+81qulWy1bKPa24AQzC
iHDF+zuu4vZM6P91pHrnmZ5Q4IrLAnmIYXXnkQpywUW3Sg4RtudzVT04TTP7TPWttkurfadpVycF
+KD35KR3OIYoKj0RlXhLkQ7Rn43fqOzKHxghWjNKZvKi+l9qrD4yR4W/NcNXIqjJYzSKxdXuEUCQ
OymBoFdQEAUyAoimVVh4o8iLVTc5biMD7nGIYmcw7fdrAEnWIG0UXixT4cqe1GmtZNuz6N7WvrHL
U5ON0eNC4e7AMdPC7sfGdAyrIueDxWaJHXC+c0XzhGwKlAeG3cGSGylZkewbiEXuxvPC8Lq2026E
kXZHMlGl8ePg6DEsjcbDQD4+hDdAsmVSfBFtfU7wGXm91+4tMgLP4LogjKwLUvrBk0AU9TiqQsYj
o5MeAgODHMai3UFzesFt18dT4fOKmkLMJoEAjwZMa/LhTs68R+i1O3gnSfnCDfBLz3/qtOA8gzMZ
JNxEzvu2NvzrGkGTu0bbovm4ESNxuQN/c3MzxGRvfwy06wy1bAmFNHTz1pgQ1/eN+OhGnvdn7DGp
6/YQwXeM0y0UUr8r9LgNajSgv8kDhjSNuRRYFgUnOL36/40YybCoMzbU2Xcg+VD3us3pjGo37Kwn
ueJVgyrA56lXB80ZYi6pLFMvYDKYRDOCxdUD5hiJDosCW0bJb3K3QsMHl9QG+QCf+uoHUCyT7H0Z
Rh1ToRiIMFkeccb0cgJZMwN63+wc8tEpFthOBWhibGy2AkrO3V0KZPirVFMwUIQnPlSy8qI7HS5L
htyVHTzwb3GiDfgQAfUcHEFrYZw4nwNUpU3OH49QauqtushO63TOePx5nnZQYWq2jwBD8LXS0PbK
wE9+gy8awLORcCHiPHo6nc+YtSGjpVhSZGqS02lKdVhxvCYOJMRjAKNBENBH6GdFeK+U5jxucKzz
vHfsXoMBWBD5tiqWLIM8jzxJcDnj95P9yWX+a7+qbexLMZwlyFklpuLHghuTFCIsISXppDyIwfK8
g6E1sf6S4Cw7T4rIT4ygADhPC+lLGH1AF5Hn943cuxBvaIlx7rgCO+K+JVh2OQyFdU4ff94CuEzN
U3H6o6/ZBlU0Mxmy3zpdTI9fhro0TJF1gLmj5wU3saLJwIea7i8mzyLZEDkYHUjlt63taKTxVWwM
eFUQTddYqikRdTEnSGaUXGNzWC06POw9aJsVvCMvlhp5Nnui709Yn1p9kAfUFF01v3Dwfib6tB6H
RrI/6iLE9cCiDbMkBcHjA6lID0WyXb2qZhLZMoZzVsd5WcaIqgMnEtnAMhQX4+KqYg5Lat/5T15+
G8ik1Ks4VlxTMP+g4eRJRswA+/94KZlcyrLt4b6VNYurEnaQxS5d/3c0PZhV3IeTwynZNJ58bYXs
k7NmM8S+PZdAga9jyYDPPYUYMIFeQH8PXiUgMpQm9ifdfmGDXlX4sGzXBs6RvZydPQihQo6gdHm/
KYWsyHdKA69d6hZ14XX88PtloMzrx6PNIvS6uXcPWIlad6KqdCBvkf9VyV6ftI1rDH2XCPvFJT9I
fAxfQh8L9Qn27PDH3+cMAOVDef5/cgk3gNTuLAU8aZ4PkFIr8225DMwiD5NRtU7GDaeQE6qPsRkv
qqw+aq8iMQV6PajR7laZzJriKooD/bahk4XAsobhMmbap3mptpspJEJ47/RpRnonp6MqbBb0sYpB
qcsgjthNr6VG6Nu4cQUnjZDxPYXUI+mpk4p5JGFkzzTl1bbnUnrROZSOUSEfnUZE0Xse+HNM37OO
wfym0tq8R22MOoTiLdBsT8tGJ5WmIsjYnyhMettyB6s88tj2bcX/lYnG/dMJyHywn3V5nDE2APJS
0d35fNTb3AmeNRsTBBCG6GZRHZswjD5IfntQj7ad0cS3LoFyKR1BbtVtqJYcMXnemlBRERyV/vwo
EX0OlkzM9O5nT7vL3nQ+gvPmxExoXdRm5OcfoOstS8q4IJn+Qghy0Mr740lMStbHmPyfnLT1oSBY
X7nByBz0IuTqMF/uYtrSvVK0CdT+lGgtxdV09q5npfXGW9t0wz77trGiwWNsiJZPGQzpaz1JdFjv
Vm6vKLvdkNVNaSYEw6236nWJ7Jvpz9isYKJ7Z7YBHow9uPRAVSrJdYQmR58Tr7qVb1g1/1tIYOHo
A/WdVwlfeNL0/e5YSOFxzEjpjFQ/rdB7UAcRAo+EKs9JyBVOAroisE7tvqcOkSz2Vu20pD5+SjuW
em0VF/JmRGX9RhEvmbjaa1NwE+M3PxsJSMLS8ggngfwqCQeXMN2+RGtI3tI63UwaotTyeiw+x797
zkfb87DDYV2EO4Sx/zU16EWt2r22waiiynaxqro+f5NjDo93jLDUiSkUKcebXOLgKVOlxtknJER0
O8wAwDYG+MOVObLKC1DrOxvwD4TxamXoP+2sse22NTx7ISVZ5RTFcAuGowhS5Us5+tvoilDhvR+z
HD1XZAl2G+Ym3PhN+S2ZZjjvvbNXxdscXO6LQ1J6uMVn89KE0kjU2elc134UJaRCbrnqlCnVq8CX
/bNkJLD99bqdtcGrmQzDxvaYUrqzJvb3F2QHazQtKBxgRpd4ygDJSqh6S2QJEqgR5CSJvxoyYAWk
rBKew5p/zF/LidFc3Sa5tjeT9BV4aMm66S+vdWJNDAolkhDKEuVDpC22DbfpmaAxqNDFkjfppbML
eyRu4U+xcUz9AbTzq2rAXOD2iSCLWw/qx3zhVmM7dW/6lU8ppU1HQI1xfWstDmwpJMOFFa9koidL
YZ4QY+0YVy/rXFi3tknv7VQDu443ibuZR2nFU7HNogkfavdz6jHXzui0pIA+Q4AlB/ZWAeG2QamA
pTmkVXqcEwyAEUGsCvx7GVmineGrdULr7O39a7/VddrB3YEeYgZxqPzmKz/OSACpf87uolXQnnkx
l4NdJJhu/CQpxfKEbGKaOUA5+IoBJ8UCIpxfwLAbnAaL9QDkBrro8Uf8udsFhUYW6phPRGnjLW8E
ERGXpI3K1CCeNxF7tN6zaYeIyJIYiNisuDCEm3s8kAZ3yU3DgOa+RKLpsmBpR6K6REQRYg0i2Qgf
o9xNV7H3ktbCefpzgn7rPSQA7RGoa007BPb523ILKvc9j14doUpevXOKZ1AumXNHPgj3wzYc7rXc
d8Ioxr59tv8VSVN7VZJA3O7j4e3dKjvxyIrOog4Ywel9aba7k5kTZRJ7jG2c+SOQF/L6ef1Q3DUA
IEFDfcw1aqsm/yOHfPh3d+j7ghvEEglHq1fGtmYcBXzswk5F9cFkJl7HOenSVgqBLMBtplY3l+J2
rvLWeZOkYiLajQwc+BDxkcnmshKNmYvKr0Kh9hwttOCmYkz9E0hgQ0aWzDOqdVmYJC1uPOjy6Btg
JHq5akK2pQLxcTS+9h00nGDA+utAvcd30ky9+yELpBrWBkFA3cRM7fO0sej32NkUbNAaN32NmPOm
D8Z+ElXwGYRZich1bx0C8yGP79zXmPBLwAskCRBQp6i9npGMccIPubyKEnd6Ie3en/tnd0AyPp+c
v4fooIz4ZMY2tQ0hqKXnSwHAAou5NA/09paTEmERoRmdgGzgXYmiFUkUVtQCpZ2doRqzt2yUxnKk
1r2FWtjee1tTB+PH+zqye+JdlKdbv6z9rfT2ZcrOMRK9nq5YENjVDNSCsGMyfRw4i6BM2IEQjTZK
w7kI8ChImrJ45J9iMjuBboPG28lH3FfMaf+EpbKKOMnx3PE/G1Ma9VLpgVVSpxzwmKNrQs/taThI
CQGc9qTqjyMY7K4AMF8P3lV3wiWq7pBNEk44FhhKRet0gWvh47WXcgtEsggNBUpm3Ofl9KbrLyLA
7XR6gWfYx0J1X15maXSlfXk2U2RBSDtMn4wpYFtUsyWJECFilK2oVcGyEW8Vwa0USH12oWnhMCLD
komMQIncFnHVW+klEwYV4i7koXRmoxf11YHexgbekSKmK6FzZX3UUheno2nOkKyWT1AJg/Ub+GI1
J2x5FmFeq1+oXrew0wwhnEDtLoIzNtzUzL0evyCJ8NPBBuvNBqXUqGkWZbdVZPiNvsExZh7lKbEs
a3nA3OnMKc2h0iuK/1Y6Wj1mGF7spO4qgE9yheKndNsbvrgJ6/ssL7nyc8EnAo/4sQyi8Doyqo6i
LSYjxl9b/+IGVx4O5MN+PZdLIEmHUKn1gBJEfU1uYp5eCb93UtDm0uwnc36f+ZW5krTmYse12IOd
sU0tsysuyHSQKmnrv5MN7Lh3SjRkta6hve1o9+XvBbymHYOL3TJiYLBHuZ9qzSbqpYZq78bd51i0
xoFQYtwXtuyJZTrz98arnhpvY29G9OQe+xr4ktTPPFLuYlq8v3KKT9254T92/4ayCf05/YGjnKjF
1EzFPVCiI3OrXoJjR0q31Is4JCJ4P7X57BQFXsHjdIajrvBeMeYjbSJGWbz5pXjaNeYrEWm9Ite/
pd5XtSRF/OcgE2/Rt733HgfSP/yDr44lmC8UQOB+GiEcQaz5yOoOCaLlwa0eJfvgBU9MctGMZ54V
/YUGIh4wvZ2RPhKSpRsfrYjgYujUaLOJgxKGmgwyXgXc72HT3iq2yQEpTypWpiDA1rhXqm0EdIIr
hXfU1oygZ2mSPzYFE4ZQrLGLTNgsnQ2lBFySCd6hmKl0/oKSB5SVY5z+TphNl9uDN83nNUr65iTL
9eCl3hGojGTpwQ1VpaiMzskQqVJs1vVYv38jHHVpr1y12qzSX+x/S9TH4SPmsgSGyX4GjrxJWmcn
N5L9kBt8xff0VCWkDDrxKNajuerP6bXqDN6jkHqP5uH1EgljgjuVpKZxvLneFTm33hQilgX5PJs4
MVvOqMm+ttig8JxWR0yJxg1UsuHI6f6zbCp747FbgRXOS2imLVL8V0Qm0DGGsvXM5iA4V4I7snNU
u28xL+9hSldyalvH1b7XF0LxFG4thnmEDeKMp9Vb2qgnp4IYmWHi780c+u9M/7FUeS7hCUYjXvgY
eL6HmDHVXqwJaw+1oFBd/xuT/3VTLMdbn3p/sZcNV1/HAKZcKrMaflRMAtqslQxdeVnH5Wfax7KR
MghQyqR48ELPphvZYo/oAqfwWNd+ZOsv7Myp8AQAsUcCSIzk2vx5n+6nfcxYYtbOcmCIWgY9ACHR
g8hu5zH8EF6BfM/+hTleNFqYayZU8MJ9IGht1NaCHKu6Bi2AuAQ4bicDYqZZ6ZH7MDrg7ulB4gzB
85hjxvh2DVJWgRgUmdaLjI2cQ7ICMIgoeoE4T2FnazNt8QVytGhO4fzW1+fLr6n1fWEH1Mdz0nqy
PNil3t8KSRbk0e/ySMNOPTb7PgsXzywPeBSprV5Avko5LAiEDf9uKushoAOkcuO5NxbO1CMOWbCz
+XtKB1aItFr84VfB7VEdoXSXGh6GbbJZe8tLtWLFOLk/sZrE43LtE1kpajMvR4eW9+wEbJYq44jN
WOPm9Osokqp83bQY0TyLfyBBBV/o6Y/V/75K1EC95OEvj5ezVKz3MyI1ySKifPnJfCm6NnObR/yD
gcwYZ4YEgMAYGD3zR9f7kteXUGeGFpRw+6sR90r2awXdzMhZM3CC9lz5hW9xx/94BH3tUhDHSdJx
f0yMI/nJ1NSinatqhQ6BVeImiVfg3lpMw2p4EFbmnnExco/tjabSzkNCH4mrkqCyMViWNS0uTMhv
gbmVNaiHNQQu+vR8ZLrXPIBmtihL/+7GwKqvTEOlzxTp/0kVyiX1UpAsj2ffTSKOnLvyyhPdoUWt
E4xNFMWXYYqj8x3pJ5auen4imVTm9Z9CE0BDpknyOwOgkchGnNEv6zUafF3aKJPdKTvOnjLX7XXX
wfRAV5HkfTuZ6cnIz7tG3p8pbfKY+pTVOpxNn9P0JKuW5RyVtGX4RdEzjtfmFn7cA4eBMlnrrnSA
nrHLaQLBJ7/G/UzOyldJU1R9eF6yxS+OSYZ5lt8v3yS3Dp8VAiqmD6T+GpnpgHYW9amDl7mwnyp/
deDM/pOPPr+gJx5uq/zK+dqGhdi87BigOVHEwRYl8pA8fwCqBtSADCBjnGbpoRPcf3O/pU9LDs7D
Pc+QfR/43owoFYn+/vUzjteOA0Y6RiXyfHQ4IT7BACYX/6HWwDPkztX6122THjqelOvNp6Lt2KH8
TTLE0biyLqWw8jLmd11a6C0GGIRnnP3U4L+GzoRn1zb6jtJSkvKYC9dJ7kcspPft8YgXs2o+3CrB
f5t7YBJK8ToHFvnqrufTIldI3LIPVhI3YTuiAHnwwaXc5xPrtbi7IhCBiMkA3GWCzCxJmF/pogkk
CEixaHc1yNoF4YX49YUjoJVgWnq6OE1g+XbV86/DyrExBGWFGdJrsNHxYK4s3wKbgyZbrxeHFl0x
AGJ/6ZKOM9/pLxTaecdrGncjLNcL1V/VsZWr1szs+pfQIU9FyRHt4r2Z+iUICz8KI2wngDviSwkw
oUyvqcQxeNSOXYzzFerjzi0BCIG4m63aE+r2gsIt5Dv8t6Zvv5n4BdZELxPXu42oRW8ByFtul1vX
Z/FJ7RbQFPjvYa729ONKyLeJxJZw/u6fK+YbM3QtESrTvnnewbwKS4vIImBHwQYWVIeYgwfQh834
LakeCX1Zif6GAZEyfxVljpnRyc17BnNrpQeRhWw0IarbhrTXZMyMnYqQx+ksBTRBwsZJ+HWbCFtN
Gcqs8KjRDfTtvKAg6NphLaU4cNqIgIJvUxRJGUQCdjfkeRIwPHUMo7inUTvD5Y3KLTDMFOK5OFhN
bjASNpPISGoR79UxM4sxUY9q5CFTF3v/L2mzotD09P5krKX5uYVJqFSKGxzOuwaBvKJygnCVZvSr
ujLsGojtyVTzxYAkS+gxwtDj7TzTG2M8V2jMaMP//sn8+8RgdgpfKpty9Mpo9MHL5+0o9JKjv/IG
ynJ1lJfwJMCDu1Lva8ssZBuzAY9nM2mDYe2eIRo19zi+0fDrRa6qES3+C/waLO+1e0XX7j+eLEEB
7vfvj1GcfURpsGInaI3UM3Rkja0AftU1M4b3QYDSFUj75+Nb9zeUpfgu3sds2MsXEZop47wWVGMo
6OfXSAzRveDVA4mORvZvXEaB0Fe+X6QvvzUWpZYitJiwG8dniNbmKgCURqTYXNwmu8d2ypXeDOHn
dDOv5ZBlE6fxSqm+MnC+qsilzxxIeAX23/ZH3jTgjXN7uXdo5jFkrGb6+Rbaskt/Bi1bAclErZae
l+njcFUZpI2YP7VfKN8owZ/HTx5LNJ/hlB3F/zH0CuDRH7WJ5SfL4iXirGuUBq0n3Z2rp6t9nvyH
Nf1WtvcrSLohDN3b0Ao9E3W/hBxj/UNH6lulF098iJUbcHyqR7Kl7P0wBGVFJjvHKZAbFM8xNwS9
lI362wGrywXm1rybrzv7Ai0bMkFFYJXcrkTQ7l5geltT4gWp5PctN6IVxREtJ0TcFuk/g7OgkkQe
Fnj4B6uxaWeX0NMtgIStHvZBG7905SD18P25E/CHWYuZfRTqwfkj4WBh54sljsK6skiyC0W3YuJ6
+Hi8imm1KQ8RQtuJc1ErZKvM/gYruuequIvzUPdW4ER8N3vQi2qSBvEgTwVYseBgjMfuHHp0xEN3
VaFYfepdViABgfqeTQ58FA+fTWNpdbjr1wZLFQH9Q2pTJVcDZw9KfCgdqiJeIwVuGkWiU8ngd8Sh
thO/81RUhLimmgaIxzp85wmj0GS/wlRaKltrDteJcOyUcH19W3oFkAI7FZSjgJBtvzVToq2JY6qD
w5HlI7wUFaRuauMVhn53dk1MVmIx/ZrT88/w9hJEeC5PG/PbDoYu/NDdZo5tyN9pqQ58XSck6+hk
wik7Gd3X/1dAeUkX8ZHMPAso3MqLHbYIZaLmexfKEpxwhQ4F3tINeQjGxDR2/URjeGP0VH4OYkL9
gtXrL9J1mx9y0uIaOIVIIMOf760PrjRgVHlttZqLVMX9kBtgEaZcZKTkzPR1yl+xznuLeGKs3S9P
md4GRqslEVrXeM2hPVpmDrb2IseNfacKcXJhADfN9waP8sO+YH3YxKoiY3d/UlxrYZk0V0wZZrwR
144saNAj+7ZsOuqFe/i3LQuXK9BvbONiLx/gtO3CmzHGtFuzQBAfAbTtABhWniJhy5hN1rgUJUFm
V4rBM2/12C3qm2t+G5yqN8BhidRXDQ8hLTn0KvFJHZ/1VfSyXExdfTPzMCpSncZAWeKwCkAq8By4
laWxCRC3MrWdbw2Xu4cxu3IduqTTyqKQoWTc6XitibL3cokZNypIsLqFRazmr1I/wYMQ02MHEnS3
P99/b1KAScwHBnt/qHezCwOxUnt2UXi4WrQ+JVxlRvoIlEk/VtDiuHopy8UpnZbL3B6Jl7/jYE7r
DH2rr+ruFVxBOY3v4AHJBRjkBs8diyl/DjgLmE9BFbQCwgHJmUb5FHWSK5CdurroffR+gqEMDV3A
fxHdn6lcdncqfgCwednJhCgxRtcmAJlMWjNvAA452Q3ZAJyaDrDn/Lu0bFCy9jFdfeoELCM9gEhH
bm8NMK30LO9b4ttzz9v9CAAT9Hzdul612hivrTk1yLhRFtErcFIXVvbjIx8qlfBg45knpTLHforA
W0tOWpLpx+yHeET7lCBd4ljn5wy0BR1IhIBQCheAVGov3InTkIklL4Trm9Rna9t3Ravw/FNL7q26
uErfpS+GyyWmkouJjqDz8gWcZXVN3fspBAVPo8MYdz4ct+ivATyROcQ2J6QJDrM8TckgaNIZZb3x
ZtNQnU84VYloAGAXILiHF1d+a1idJVMWe6EIDvHEVC6vOwJWktdkgA8RzNextb4v4I5IjAiXX3c/
rcLVuv6TMMrx1FJA1ngVOu6tbJ4f4A+2DJ1i4Eu3uwCjdr3ZvM6URri9eVITjw1zb9w1POIad5v8
6PS77qV3rojxCmJFtlK8HHlHzvZRycJrXHWlCBU846exRve24UwuUQjTsIA5uyScu0gMRePZLliB
ddkroBVzEZNpa+NKIo0I7Atn6h+vXNB5w8D0cHlja46roNT0Wn7AZcPETizDyihjoJXf2LJhCtKI
djjE8a/XrKuq0acY/tQFhJwyGO32pj/4LfJpvOztiGSihPc+XD8uiAIfSjOgVBxrvggUlmFLczgb
8P9Tqr9E/mIzMtgF3sC2FLGXu+dGV4XVGp7JKXP6qQdDiA22jW+xLdrukL3p4Z2W/vfdfFYas3td
AS9MVvPM4rI0mxUF2An2wJHFg/XXtG8NTTRyEG5AWBGUtgaJukPHmXQP/hI2DOt7JHBRlR4UYWEx
/t55sNG8MlhQfJYs1poOLiT+MIovwb1kFkBMpx6obNw2qA+Mm5/ysaB5zo/0/E/3dNyjwGSD7dbr
a3He6kDl7XSlP6lp9OeXw0nvHKDBr7X+iiaIMyDS7yALXk1bBu2hk1dfFGnmw2sGKiv/4BJ0UkC2
iGDbP0WFFEn5twM6pVArovvPfgbKI1yKq/wlBrGYiEMacrVqB2lLyI6MxLSumBkyvxNCZown2hTz
LS+TS97KBHpv9P4hdzdT1fyOKLbSHXC1ZDJXZm/XDc6RlTfK7Mk1pmQCRzKqnvhNPyJnMRpSv/x3
hIFi97iKB71aYS37GJ0jCITr2MAi6fHaX8N9F6J2Ha22iPpIbMBCRJ2IN0JcUSGXCGaY9x0EvnOZ
MRgH/UbaG/QtHY4yymTjfENDBv3piOkvCNNHkCqQzOZE+BbDQKn6NWwm0ghNNKnh/EykD7kiISHt
eeiIVC7IXJJHvQMocq9AKrwtVzVQxJHUpgXSh15h6UntNgJrTYXaET6civW11uTWqGMUHaG01ZId
ob5KhgAC6IyxP+LczCvhQS6tvq6CBB1wtbj0Irf77v0xt7bCdAqIyS8yN60m8KBvb16slY1IjUs0
nzLYLG6jWigl4stgnsP0pjbZsFnHuG+/D0UWP6NeOYbn2fDqsMl9voq93lz+66ua/M1+K94MJWwi
SlwbQiohNzzhPZuVJYZD0cXEBh3ZZCQmkLs5gqT+oXin0w+SzFTTH0A3aaZ2PI6uCfN3RaP2X2Cp
cH/8eCDwiEXmgRY0mSmrPOAKwO2sKYEZL/Sx3VWKdIo/lzqD6BXoxHCeHHTBI1xkbH964bzrNjmH
muYEMz3rAqxpSbM+WgscidRygT2fuQKx3hHLlEwdJyCC6MR1S3XvqG8hTMcqvQqSbFr/HE5XQHxJ
wOtEziw15PeKis+f+IEvpCKMKxXmJsE9jJFJVsLftHULS3DtJX2SIXodAAWLyxo9uU5ECxqLHtO+
3qmAvUhJpBiGdtSXIQLK3WKKXSeyFtkYRDFUzTO67rGdjpk6eelrBvmIaGoSXPGIgOMVMtjomP1a
b+lWDHnNpu5SOzdSU5EyVJ+sESc28lTfRFWS8YSj90+/F8Mqgt7Sr2nUjZ2sxdWXXCEdWbaGCXHl
xK8kxnDr/21KIQruPSYQMMUSfXkZfb7g0KO9Ju0YEk/CW7Krnbe0fjnHFpP7ezy3nBOM0d6ChjOy
CAFmRMmEnaee+xBWR4FYl07pNbae1PeJ/dYmDOpDHPiDwmZ74+QrgEqbenIfDN/uY9p4+Lu5BaPY
jyftjW8BR61CbuUZfqWXevOoY/g5p2xKJl8iZVjtOh1nO5FTb39Uj80SQFpflH3ho696m/NSpGhh
JPJG10fLYTq9kwRAuMa4jinsqyJ6FMaJoTj6uRFoGuaPaYVbn+gfeIjds3z129oVMNfH6i/MCaRL
VvE5P8AWaosF2UAopTkshxt40CJMVnKyjgJC4ijtYe7a+jXW87oYfhkCEUEyMtE7rUBiu6v8WlQ8
h1l+1ifZHP3uY8RLmRQnbiGPmp6K8N+eY4Y5rYIROGVKX0wqFW4OV/+LYcc8+OFz9M3NAbyZhP50
WOv2Cv4+4f+uY3OXgYz9vSCE5sAb25HKW8OTGgsUlH40258ai01jR9UGwei1Zs4p1acmVxK/LZLG
yQgqmnDl6xX0pwrkn9NuO+GBb/v/uj8KHecZcEsxjDsgBXRkwOLvl52V2+CjeqSs8w6GZZVSWOEc
gIXwex3ysZ8apSooBNO+dYV73jgiT+Dfvko4tWhKDXqizqF8ubIpZkwG2JzyB7BtVAoiJfqWoA23
lynUX6RXjEheTCBS0o00hrLsXNY0rZa8uAh3wOUITX0+Z7jQK/F+XvsqBOFOjTx6d3WbOi66JnW5
eDgElOcpP8jx45NUH9nxTwSEIuGnfAacnV28KmVqjnI3brVM9miXoqftmw7lNHKWNO3VlOvlzZvq
Am3sOeA+JjbNH8B7sZgRpp3VkS/TN8kr8JpbQfDJdwSYCloSZcNUM6fDrjExuyFXiTvfnpSuBGRj
YZTejSEvdlArVKYOu2ujNRRhvKBCi1OxpTOFI2+gIGr9NwPNAoVnP6123cLC2E571zntX2xeTFs1
oEzhxucj58NVF4lkRQYPfo1pYGTgeGVJbJIcr630dVNTu7LJ47ooVbKC3HD0QEaUe+0YwpwPpeg9
xYzyhQcnSmRmfpmAsOgAHDDbZRUfKZF/d8Xjy42VD6Cchyg9c/WtoGwoT6EtBMWWiQLlfXhDoZPY
gR4xhRfyZ6UuhQnIShf67kEQSVabQVfZg7VINX7Z6Bt0QOV31J1QDv7XVMh4KS3LvRxK0G7pS+nr
ZptHDdXeb7rE6nActIXjzQaLmrCFSLbMOGokQP8gBzlMCTkJzOb1D4VjxIhcAXWcE25MxXw5VF+W
S18Y8Pgcrwjkox7HA9rfFJyPclCx1OR38tGuuYERQPlPMYP0vrbn8JIrI5jBI6yIIhR21nqaEtei
McuG0O7zj+qgunfAYn6J1tSDP9W8d21wqXVOwWSP8yj/0OSmkt3hPBtfHbdpGo4nlXJwjm1NHt02
AUbJdGZ48DbS887gm1U/UdBRBke/b8iyqINn5xQPjFc/dN55J71y+WpvKqgl6DECyCtlL8Nq818/
ByfNY6IT4UccyNvjZ6voh2ndgSCiIMQ762ZNhZ5wuKe0A5X4zTkOpnz4jnqo7Z4QOjEnlZ6hVk1k
oq1cXdHeuwZWpw4z3jwKm04cpC6qPwiMSn2pYHjnPJStii0sa/P64AQTgwqFikoE1ImS/PtIFOEh
85V0n5S/muLWm7Few+a980wZK5L92pA0VKwBNwAJyO9PFhP/5KtgrDJk91pMGIH16di7NavBmvRP
5i6qcfhYkGw8fWGOdmqH8Y3RZQzOqEcoDkhWKzLvuEEOzBHAuj/iNr9MxgXvHKDEXNYUh5qAsy6d
XIiFb6kHD8AXGmuDj7yX88K/xwZX9BwzpojO7NUbqU+LLy7HJvRzqvsLtHyKUNjZZjSdRjZL/dUn
U/DoroklF9E5scCnbWCYrox3/C+U4mypIqmxf4H+G9V16u4mWk/WXOnamiIdWNWcTGk6+S0FHY2N
ijNYlDVgrBWRiAL4x+gXVeVP1vKPA2GLqSXXbnavttbdYgarpEnlbQMQjsbrhFwQCWPJL2Ru9EP9
RCbC71mH2Im3bGz8Dep+QZZaJi909d4aqbwpIZqEM8bby6YYOEuXeYcKP0B8+KNDqtEMjMOROG92
RKQAwuMe0J8P3esAMfwVSjyQRihMM65PT+IF536f7SAOFpURw9GPy9FNJH1+ltr757QU5x42JK7j
J+yYnh8RFjur2uoVHObgtgAs867GAOm9gSxv/qMgWD0RLVNLHwnIFJzVnybQfWWWdaOEw7qqp7nk
exrj/ah0+Dq+e/NG87OGTi+oKFdgAJ4BpAFQXkuGeFunxGjC46XerRqH+KD2q8Q1RJ+1LSwscS7W
xNRcwgJsBpdhYAr6XQPuPtUlLPbpHUnaOvBFOO5MQ/JZnDxR8Xt9JYMzh5QaysRgufyurZRFX6ZI
K4uJfVWoOlyZKFxyMirEktMRIPLiomYdEfHij3QDADqNri1tsPzXAn5/WCX4oel5svGFOY5TBETQ
6dIn2DjKEMijxO3FV5mtW4oiPvjke4cV9Vl0m8nP//SxlPx6axHFdjXNHcIapoABglrV5pS873k4
FXkbFJx5nzU6ajdgF6kTmGoLUOhRixLSQ3yl379O5PyjPsPaTNKcg9sY1xnDpF8+s4IONW0wQGA7
yi3M3HrYBQ3CyUg/y8QztoXRT5CLBjOhl44qEksFfYLYO79iQ7NpbKvn2DyodSiNsBVhenKw1i4m
rHdBXPlO+6hrg+u9Bhc6Y+vpt4q3KicfCnGNzb65LTT96msO98myyoj+YK3CaLxsax968FprkgFK
lHgXQp2WoKZCa7WC/Tmt6TnPbrpfDTlRVJAnf2QZfvnavorTBFS8UMqFoti3WnaEttr7o4jd7hM5
7yidX0kFvbw5xxuzqcufTjhTvUkdL/3YrU+cGZ4TB8gY5GpdS+uKaO73RWwwx/HJTJ7/GsHw+fQQ
iIErEYCHv+2fcAMbCQ5hAT7v4n7xcZJy8gmjBpPH/dJORjwhdXVbOATmmDdmS6gOy3XlIUw0Xsfx
XC4wHVJcY0Ru0Wm82ZdRYyHZeK25oncH+I2cQjg/7PlQCiyg60OCroEVjrKhjtJagNyjJ38j9hBC
qVwiOw/geLorN2MGIcN2LLGXXqcEGZPuWVLZj/fybntjyxgz9lqjJvm/xu7SrtwrIIhTJUqmE1we
IN5bKZrl3sC/tLl4VwFrHYeS3cHf31JUZhWcXwdycN0QzdfWpqkvbpVYMG2mFpsNNPZ0EY91N79T
3wdS1OE5QuSaEFDfD3bC62Pfaz66IfywCopqsSl4E1pqxJHRCqmzNs55JZk2UCgPluOGDIWOzFM3
9f6p3+YmBUkPL2d3wbGPwEdT0KtoYdU3qZUqGXDZGHf1eJhjdySKj08hoDfmPUxApAUqL00S6miJ
GOa8DgF6/YSc/kAU/PX1mPLOG9mvQrKyqoFhGWkMvAFEoTqadi0jCc/JXGOCTUte97jgeS95ZbzL
dKGzE2vTubME6OXf0P6HPK1kRWUrnDk4YLyCQc1YF5xVQ2w4+0kGWF85XydyTUiD8zX+JkE4INJx
ZDw7adWgcLLWA6mJ9d+qLMVTsHvtzIPZSvsR7fVhrdanJ/wA7bDnL4nZrapKi/2TIna6adO7AKzd
YwH4MJvry3YHOugSXLCMzOLCt9oEVkB7ybMuN1C8sEYD8ZMRBm4f6G2Bfkwq0P2zzTqEnij4wQNg
fRai8JRrforuhN4vhtxgvr070k8T1HaqZdpAty4S5y7pkoSJsByorAM/NahharDyPjm2GkCzDw+n
AMmPOfp3WRgKkGgSwLaPjtuFbLxENEvxsM/RWrmd/uDI+0qguiJIciqfCyZWKq8SbHXqZ0b15twC
DHzKOu/6DPcq5MnoMGYAzafCpMTOp4p8u4wijQrbBd9iEk+iTAJGvoqrokhztxm2IBkJwTc0NwcH
4kL7qUv+VNZ5LjmdoLnqcG7/VV9yb60kzxPJtiHvHL97zd/mDTCEQXluvmsxgBZlLCpmrbtx3t7/
BBKC2uIokvIRKp6EHydxck6PMUkIQQoujpZ9mhE8BPZvHepXKz3e4dP05npNXA3YabCBUtkzj8Iv
JjqHS0ehz0tqwncPk5MPSfJFY4Cr+f7XkOofMqO4e2Qt7ng9kDa5P9qkgVhsoU468PZOdIgIqld4
k42HlvbO5RPTg3cQf4NPbm5iPxY+mIVQqjlzUcEERpcMfQ6pqWT/c1BEzVgJgcJEpd2LvcbRauUo
07uL4EZx3TafI446xlAG0UGQtA9bt36HVLAhvfeNVIjmfNbtSyr7fmMw5HeQgZFapZm9yyg5hxwM
4qYQVH8oO1kZleI7sj/tW26IEJfFEKzHz8OttSJbAzHxli3rVVWcozFtVsW5Qh6YKx2kTgOqSNQJ
BBPH29WCD8XrmAPamGtcRkksxIX0ZY2NKg4NFo3WfAOwzF10UO/ETVjBCA5niuWDGBEUI9HLJWjE
J4mxaHBHdN8FOnwHQUv5XVyRstxm2qtH4pH6YFw43ZZkuNbMWelvP5/iEtCuy621ethetOuSQ8gd
h/tK29vg1xu9UmQ0fbmbN5ygb+TRlDLLtEAS1LbmpLc07r9NDlftuI8KJz5feN+ywKNnW/X97VFj
g9NmAm4hEtYZYg25TkIHac4uoSJsbhyN+hAguz0JwXgPukGG/mpCq7yQ2EFS46Nyfn7uQB4R5HDp
CaifNe/U6LW/LzcFIUFgdemJEtpqH4EbgaddLq/oG81Sq4WbKayrtwPy6JSbthB1yAqs8pcbD8J6
KtsgDDR/R+sdOK74j2dn8TnCfAcvgSRS5879F8XLfeR1wKW0vYqW34XkRIW2NpJhghCVHNP+VZ5y
VZZJt1Vqu5w3SW+rNdwGjxRfTBr01zCUJl7qsRSb3mvfeOD6RgBXG4sSKXrsjAqfmO2+7tGaQzf2
a8/sKlD/ZjMiSsVLc3huSvMKHzBWSwRRpQHvIcIgaEPboQxgWv/319fF5uhti55cDwcLRYVqfIdS
hITRfPP82vaCQnomM3YatszugoJBF9iN8wCmM6qa/6qsXH+mjewu+9gn47wBpNalPTNpw9kOQry5
hetgVv8JqRFHZm6MJSJBZq+57v1kJogFFIZRaSRknUjoe0s9VE9/i/x4a6O9ygGUd45pH2ZRSB2A
grfb8VXQ/3jaz+KHcowDKkBEBwHWYnbglOrbYup1BwJcnT8/Sq/6/jfAV9s5x3xJqSI59Rbcur26
kOKilacHLgeOgdO/mjIGdrK3laZAf+qKtgRr5vijhpXH9h1axVYj/Vk4QYifo3eHiXSE9WDOdiRM
cHyA8c+4405DOijeNHUKAjtSWyNrbdU8zdWWy73tkPLOF3xk/DLoYdAXFfGMKIQnFow9EPK1d1o6
GMIkGqjj5WuHW0VckKfXiq+Wkdh7z0NjHZw1i/DdksczHUkBYXA4vmz7My4+A01IYUf3JVPGHOeK
BsYan4RzR+7GmJ4sW0R0WE0SKhmnhIymvUnLlSzNo9KvoaxFyNpdfFMlveFlA9MKCqYH/rN/HKVp
8htT53dW4y+wsc/SlAhM7P83adPsl4tnA9j+kBp4+z6gMwZ2CJv6gKiLj1KgVUZieO47jKdlptcR
lYwrK6P3esUny/kjOZ8Eo09uKIQkEPfw8oa8orV65fUcXQcDPPAM10w4NSqdJjZIQ7W2YSppvE8F
xXJ1w8Mk3jiuxLoLYm+2k1S5NEIj0Nc31x21zsBmgEIr6NCBFk/3ACQ9umNKwA45c/u115Wx4J0D
u9/ic7f0Hl4bpwm1a40j6FOQzUFrRB30h0GVEyJjt4oM9HCHwBgc8m+HJGrUJABVom2BSRcvGyQx
AcY5mkTCIZsySt2R2V7N3s72pGdmfKHHdx4NhD7dwroFR3ZbY5oisOkv4jbdPXu7KfMOOzBS/gD3
lX4w48UTIvJ0al4bbxLFCOjpTGJxO2uaagvFlWNeOvBK/xJ5k3tg6juHs5U0kWaW4H8+qxyoHf2l
9S4ndWJicInkGx5WHm5Hm2ehTTZLLZnwTnIcND6z17I75YI2ux9loBbzVf4Mg48nEReGm2p4LYHi
swxOGFruoNyq1enAQiJ/VOx8M6+kiuEECzP+f7Kk36x0qSBxXL/N7nSxZ365pai6K95wvtV0yR7Z
XfvQF5vlMKsEwOn1D1EOzx2cqxizu77j4/wxnQr4Ykg0cW5SNQCwZcNrldxPU8r09Xm1zHqvAp+9
7UFABqxWDONZRFe8Mq+jK3fQZAOZewf7p5LGYcGqwdhpryKa+UNPgd944UZytH15EfodNKNEjGjM
of2oCLNFcsJAA5SKTybfJBqjsPQ4KdBcEgEc/dGG8kaCI3gA5GbU5mlN7+3SOqY8pXgGVtz3JvPV
0CGhcp6DWMD5qiucBOq/BiCW4CblljobcMstzOSk5bEVDIA+7xRMg5lQEWfIiAO8Uwzx+nWXY1VX
WFHe66HiE+52MfxrVC7BF/Fsl9sdDTweWTAMus0DAWG7JfuMHCzJE8xO3AFIUNitwiKhXqSey13k
uLthMWVK1T72ceTJ7fyzc1j38GYo30xEVF+5ewW/8Wz+QWcaKX23wxkQaDqbyALpcs+r8mxQDwAs
eAXHzMFNzikS52HY/j6zNWNx66YuazQAsZGoyETUUCLVqYiy4qxGx6ymwsMELQ4//Qg4XSpBtiAf
rdQCmq3qBZvkuFenASZhj4uPhmSKqga+Hf122lCGU/te7D9erKLm6dfzC7Y0aSKQexhb/I8JShPW
ddaVG7lsd+TRYKyRokBstAgRXykxKtsNDfH7YJpPEzbMLHqqMEcr73FmJaXkM6qrTS4SZFhHpDva
hDaS8eUo1tvb1azC9Hmz7JUiamTg7TRapxwrxiMjF9Cbf+bgVBS/wU43uvWBffRW1pElXRs51QWb
BthYB2hO+GO1o59pJjkBwoFc4lEfgSDYyp7Jy8mCHssJoWBYH/eHoJLcpWnYkWPXxEXCCSVSpj6n
+eEoblE7REdY5PH/e3rcFkV+4kzGKJgIYobktKq6OhCpiOZCLyaRIH08czm8WbjB3R8/RMUbQqsW
ao0M+zvTp/Pg7vYeSgkrqX1x+jxlcp4ZEtwV0fv8KMxjICYu83CxfBen4d5sySS5bmjAM/2mh5qC
3d6m3xZMyw78EVxl/gRiIeE/AODGD8KFX4kb5AluBv9rArucDd0diBdLBpdnPwhuXxlxgmm5MfFB
dY9EIjuZgxfVv9Tt66epXwjm021bxLZ1mYJg6ZA7Znf0gL8p9LH3dlG2g6Gb/z1ivCBZVIUlGE18
jIBceAsNHhWgNSXGpyrIuysDHnBc+L9gWNn5wGTbFvE5iVc7ruS/AUjyP9nGOSLtKAfcbnffLpIL
H7b2QYighXCVDYNgg3uTRuyN4ulr5c+2j9ArOkIYkSQzb/oDfmem0cR4d6pXsIERhDrktdbq0oMR
2ZpKo7G22lyKUibEAPtAGMN8jA73FY4c3tZYgPICeHxMw6/eohWrH3hBTw83Ii1SXu+oLq9TksSj
EWw3rFg7N0/ASONjeRWb7K7XNMM/t6O7EgT09hVHMuZBUIBYHdfiExHfUheiE2lwKHlcpz8inI7m
sf2Qywc5eJBldFsrqpVMrsa7Juc8QqY/Myc9iwjk+p39TfPk+uUPXknfncFQJEf8y5VX9oHsTVW2
2Nl3yAbEQy0DYF9GEzBouMSStKkRwIHV0v9Xh+fPA3QRO264LsUP0t/si2P8eiDgnOsxfuSv8tGj
ACK+u3v/QVtly0chUtpbygw4CrQsZgVUQ3xKbC7ReRHlUuC34rtVpKlLK3B6J01Lu/NxoiY4AhVk
EIhHlGT7DS7arIdGMTBFOCphILoHUGXHuQbXyaSjYmSqzeJDYmyDR6310AELGjP83nYEpRye+oFh
ZeZEROtNE+WDenzGj0YB+in7kvMDVrfhzNiNMaWJxz0LRauhys+fIl+ujZn0y4CiHlgCE4jqhV/v
/zFZoP/yH0hNSncsj+xlMEa9dtN0yopHUHUCZRSVgiep6MQEp6GsX+oSOsoyb8tfVyseLz2s830T
iHYF8getmRqMyMGLaUjbUO/6wK/4TnQUdTvaTX5LOKeFukK55kOEPLGxbNjTFN/kDWYxsNG3jeRu
wtFCRo9ekdsdUMaGyGaGWCMNwglq1QA2ibJVLnKAsQrytNJlXG1UESqyxa/jkRPk+W2pXZKnXV+q
0X88+R4PgAHuCsJgzyPcwnxeqw74GA7T0ZVkQqVuIjp7GwYpdyJ+fT2EAF9jsb4wTvli3oTwRZJ+
v/pUPHDWolhMqIh710e5iq/Nl3hA6vMqHZSdREHoZQzkPzrWolrsJYyzvOW6Pbn0cOJwA3IZ/LS9
BnTvy/V/va+Mw9KvBCE9DUgv/QvEZ4KxFmiHvB43/0YzUXQTFDHxs2B+Yby+gixfCE0tXDkZR98U
+DaG6CgwQl0jdIs6L2q0+d2Xan+c67LCX5cNGCphdOALMYMjkUXDNfPkRC+b371efgc0zI4W+Sgh
zV5tigw2wc8mTrU1xHZmwJ2xhU5XFrMAzzPAgLyFsuAAY5WC0PlNykGBupSOQABhb5i6jFvSn+Dz
4m/59XK+3YkqulpG3Vo03KpxB7uSaOyGWwImnEedOwkWWkwIGcpMvysN2rH41aWSK4jvF6VlN+at
aGMJz0Yv4ZO4MerM9ItPmqeXN/XlRPKHZLVkEk3hPQ23aU8Lx/KFmeyxMuZuPY1Xxm/r7LQc5VlN
9pTyDC3NFR5UgW1KAKOjGULFzHciJaZcPvrxv1ZDBEbp9itm6+L0P9zONB7YPAu95m9kXsbC5PXU
lye5y0gYM20Og6SB5pM2p7h8X7otZzcWSGMxKhMblrngETJwZnPvKOaqa+Y+y3Q2mb/bgL9FbOfE
ziocrEHun5RW59uWn9wrOePt8BePN+Wl5tB9AQW1gF6uOQXzAV56vki2IN+JftQ2fiJ27cQe/OT5
GVS8MGMtzxZcGqU2NirScZc31Ya0k7BWvX/5PMKj7ucmo24kcVM9HRKYTQ7Z3iSLZ8zSigM47POI
gijl6m+hXcynSBiiNs3OJES6QhlZ/WoyseTW8h5SB0tctUlweuWNepb4GFcNbCVPoi0ru7xidtOz
Mbc7zkSzdmuMUbV0CO7qjVNzv35kTUQX7Cr9N2wHDeMF1OrhsIi5Odvi7shbqnLMO7+M9GzHcZC7
1MYUmg85TnBVxpZvpikithfgwgxqs62Ugtz8mEJZ0cXHbmPrRGpT3/1wanUR4+h5d3bcQhRpju3E
afI0CPYtAAq35fHjWE0M3EBHeJ0p5qk1COzy+hY2o4PUBQmvMHKHjSH9G6GlnOgaPkMMS/wMERMd
8UyrKPGgKA3Te74eudhqi7BOmRiuQdA1DRAiaiY/w24Bw+Pi4Hosr+LF0V5YUpEqCfYl1Ml9ot85
E8EBzNQsxKy2ZMZFoDAqct4YGcky7CIPYz2l2FcZpsxxKWzZ7FrAF35jeIhPUlvWXElUhW1FsjIc
fMrHJwmQX6gU05I9Sj8vGeFpBMsbEo3lqd6sR52seQE+smF1A7XUo1H0+BkkyzKVhIeHtYpR9he5
SUsIKn6PONDoGpcccOYH6zb4EZQaZcjdhYIXMAOoTHn0kPYxHyYj7+kpjITe/haImcDkSNg7UpnC
2V5L3Yv25VXcj68vGqxX0LDQUGLcEddg3Z6qZYwJ1I1oZHfl4evrDsZMFv8azLan7qYyXZLGA7jh
ry7vIC9l8lQjtH1ETRgp8WBgEd3yiIqNyKurWdSVeV+J1BZqTtTpVk04RWTerFlx0FdEL4s5+95o
hHcQcgrIQZk6ffSWm7GI6lslN6ZURDhB7Eq1TlOzlQKSEfy9T6gJmkYfXq9RHzm40dWnG9AxAbHh
PZulGjo+DKaEs8p/3kbFtDnXLJ9ngR0dT9jkyWovshiErMG5ZZdEvqu3HJEOw2YqlK+VRDUHZkxb
6W+BNjXbcEVifyJ1pWcgctqvhhN3ge6Epbu7KtdiqzCzQsptL2k00yiJbleNGUccw/s21Or7CWud
J3WbdbN72QGEPgRNoPvluzSkwuYA0WXq0NWqgSqGdoeq1G66ZqDIgYSQI4JeEmzm94u9iiAENtjW
TQEcJdz9G+zPw0jq7xE5AyT6DjXx6D11Vp7UbcZ4lJJ6Jea35g2vv77s8+cW33Y5dLG37UFasrN2
0B1e7UEDraRHB301McdpuJYeyZ566nR9jWKrZLg9wJiWBBmT4KJyu+uL9SdivJMAqr5vCOvfh0Ts
38mthKZvUF9CI3eyrllbbzQoOrmeOsCUP+Ha+C2S2+u9s1rdNrZfwURScFrCKdqnxzT39R+ciKtE
Az+/1MKcVPU8i4FvhdJvin8i9JDEM9MOvNvyDnPoUG4IbOv7pJCVQNQqDCgkcPb/qA5DB+YMuApw
zUrAMseHnfAPf+p15JQhwQIVrWs8ZqU1LJDUSXyn83yK9MDHG8brhw1FhrUi+X1eqzNgzPjWaCBW
k4Xk/O/8eiCq/3S/HL/PpAQQti6V5rcX9oa6LzGFmjHV/WYrtxDRBMYUbW3VCW7A3BwbDgyNOfSK
8kyKP8zjLtrTYd4l2HJzSytLo5mmynHBVKr+LmsUyv+7JfwaXMjBhLwRyRrZYE2sHJQEoGlLxgz7
LuMO0C/5eNNaz80/UbcbIjG/AAaDRYq8z7nU6Co0dZry57ODlNmPnm2arhGUP0CJbMj06q+16LI/
FdfwbdL5TXtAni+S2vwLdwfdbQH0UKqZLsmBXwgH07gSvRZExzP910HcKCOinwD0jJglczYLVJV0
6nyFfMzugrPs1BiYIqjHyDfjtJi5ut7FmY7yH+FRa8ohYytn7ylBzJX7Zv6YfdysfoYrCRuxx9U8
NC4O/Y6zg2dz40FP9D+TrVd8ApfVakwuBDkRQ4fvusFcXDTqH/BsEXRiAilo4R4wiQxxqa7+Dqyu
R1OLscaqGYbaD5O0K1xnduL0tIBjb6o35N69rngEsb1dqbEZudUjzLm3wVbXbmOAqSSmZ02/nrgG
MPVdZ5EddgCMy0Dl19anzWjJdwpyylzMmBNzxq+rKUW9nBu/yfJC5u9C/USMqr5QPzRDJ8MX2VEY
wtEewAt2QbVld3BS9CYR0/s7D4BHgNtBzEetmO1QKnUtr74RGZy+PstpGSPQoZzTh26QzS5188AP
emoNIA28E382LOZGlS0QHHtlqVT9z68kDn+hACaVcXS7YnK9mo23yTNqpki4yQmNralI7uF0V1Ct
8AmPp8pnhjSMVnJe165GZoo7lx8/RRgHi+C6L3C9Yp5UVaTheGpv5dxgJTXrgSAKTpvSBqx6Y6kz
FA1/i+TU6bIVXpQ67/ONxnNJJXykR1uJlSVakjZVh1DHyZyitfK3yYx6P+pRvZZGcVpSAjOgzidj
7mmUehphS2yi9eaWS2N9vnYdUfhIWHQFdg2WJQ7jBZ6kmmUHKWsdMXj3xESJlt68DK5rObtjjXps
F2NCxXdxTHUs941U+ud4JejTsoOPB0ACe85pGTui6KjoPQNZLm1dfCh+83aunZjNUAjUhuWk9AMm
GRcNW/Dtn3GBQ3wjqbSG/58msdrg8k+6BviK/k268XbrQ6F3hrqqorssUWius6u/gIUJXGIcPCcK
Lg4mtydNT3vvrbz7JfcAGVgaqKxX5vDh9q7lhZoXrrnYHy7hbaLQBkgFU0eA2K8cY/KnWfH06FZm
vYQYuOyUKUtNEIYsAIqno3thdMFQGPBQnOeeQDB5nw34PrqI2zcNLqf5BNYoxqKTJLpwkTO7LH7K
kGpTXUGE35VWVGgnWVwimkWbIVvDAoGC9US3FVDPJk6VhUtDpxAPGEqcjgBY4LxrValcEwlicLiB
7J8QiXTosqDbFI7Rr36GuBEXQ/Q+yJfybDj60YVg/U+40VYllhEblIBVvNpgYQ4TwzUgkt8Wvvk0
jTil1G/z3OxeRG3KuG37j3Ma98sqMwEbg4rW7MbazL3DgfdxcAjA9WlxFXMCIUivzCXcDkOz8QiJ
XNVUW29PykZqpzdhLI9OXDYiEVzXqBeYEjrmIkRR7wCL6W8lZvqReAUUT22xilFKA1pPE4pB11H1
j12PBmx1gNnXXwWuw2w9Dj6Vt9admVSBMeKXkrbBHqUV6chDQwss20jP8dDt6GNkvGyA/ZXJl/Mc
6otwGNoubYIETm9sDr7HZoSuADdZaba1sRqNnM33dZJqW/rgnAQETvba5+M7j2q5Ymtv+yWSNrm+
NWx3Wx0z2fv1JB3xjI5g6M5NvxrdhbYaXrqZj0Tc8o29NUbcYZBfbYvYcx56X253Nm+VA1mz1qzu
95BVPmnJYnuPW3WL6uWyaa2/7FT4yhtFa1n6UpS6ZpmAv62lWWcYzwpjNB+dLpAIxuT5NvGE+s0Z
5kLEABy+JhqgW8JiHjKUMJsgD6HbccYCrE8YxmNEIfpaVPlS66wzhFw1+ACH0ihIIc9p8L45VBZ/
MnbhqPYh+lf/awKSjlu/APJYPVsiyDpLat3BEIaI41wPek2QdvhwjjqOk4t0q6jpEzvBu6ME+Auk
/ho7IqkQuAJqOqC8/CC2qG1Sc1yFWiv6wE41L28jMedQZyPL98rY2nYAH/K0Xo8f+KGSUMs4s37+
Z1Gk0ZOEDkGk7ObtUlKcLRe+hY3LSyhiyoWNxsZquguhi5ODHGmUh6oLllHQoqj3y/wvXRa+R81J
ElGSnE4y9qZ7276R5L9YY8U6C+j7STd8ylIr88qAFZA1YgTTINcvP8cV/rq6CHc8JA0pDXHzEMW8
+jrHxZ89pVZGdShnIvcqOxKad3u0GRIXGu06kZ0pU4vCCr/dyCeLJsXyFZlGD2z1ECU6Fmlj3VG0
edkeCjcNRipVJEd4gDQaTDe6ObEG9i+mua8SWtvKFLNx7H8r9k+MOuKl5JaKXQlgKnZWL/hKdC7o
i+ZgPEXh0T7MldQ37s1ItTJNMCpoYnWx7F3tp7528x7K5i4wvkZ5+QzeOae7A7/873IPavBaKwxp
P7QieF0VuAWW7cJV4NkY+QBCcFkBEZ125oS9+yX50R3LRGhSM/arP1MffTO5qRtt5uxu67Wr1Dd5
mEJppIRKUKvJzaxQ2uYLWkc1+ZIk2NGkwbKxWraDT5AJSwNhTNCVKhvzWkuju5B/FyPOSO+GzIJP
xLERxCyibkF0JxwMdulaTpDWdXw6NMn5fpKPUAzKnx5h3IY2FVqgKKFMs6tmY/kLqjcrCWaJSbWS
oChqg9VECEpxVqk/jSBAUMa5T88ceNGg8LmKSBvuglh7oUy+Bpaq/Rt6AwOY0u2GpV8e9jYwBKWT
NkTHYpk5CvuhG/Bof3boXuZWEjn3UmSkSqM03xvTmjbeem/NM+jO74chcw31cTU/chj1RU1DPqRl
zHbjpY6ItZb4mc5PMowz3OWfKmCYNfm6LKov9tTbSsGO/DiyCMtyn4UAH8bk0qJuXUBkCvWhOar6
NiRt01+1Wh5jE+p9SfGmmlteE8bojazQeBdW8WyhcA7Oaqtjy0Z2l3mQYixWUjRYr6L1kDTLEtcc
PmbCsHq3gaCwVUyYzdcK3sB/qapRtkcPqfkgvErGAoUziXrwjcT4EjmiqJBEKfaJIC/5ryFlae6H
sLf5YvT2WTe2PhaiihGDQbZ7FprLbhBsVvHPf1NXBa9fDBwnlEtA7o5af7q4+45FVJEUJK1YNWnQ
AgshhgRkAkZ5kFvqEwuhEwQmhViqIXoWk/cDxfiqJ63NL3EIIT52fefMmS/G1y3xU/j0K1iABluf
DljA64rNRqBPVgGtzddtWHUPHTSL385PUWbkAWs9sbgrgqMzAwv+t2djv+Uo8kK4AuKsxw7vgHIb
tDTBqUh+del6M4SChsmGv3mczhyZ8QdPBHHhdmDwFjme8Ys5trzlb4XWG4D5GX3pFWLyOAYKRxzW
TdBSI7Zr1cKa5OsegDZwB2QjgdWB2fH5LohlWrm9umQ0fhgEGZVCDvUoUx1GDJRP+YuFw4hT2dx4
slddN7mMIaMKcunhHX9Je36M/vkzbC1R1eyHkQnqSqatXiD7jsl6+OeTY+tHdsc2+3SkRCO46uFy
nLAKbWL7bXn5Vawt/zniO3yqfY+IijFAmaIQZGJ5iufpE9tYUTmgaUVqs9TlUHYFEwU9aYjQZqS/
H36sX51li+FWNm6khrqFXTqu7WqChNN0a+lk8Ox7+gkl3lCsi7Zi8xj12LQPC6PZiILnnNoUdujk
ZRdHer9UnLOfBCvp3dw7jmohRMa65ZZTE9dohlJdE8qYXn3XwwY7h+rnnLctD3Dj4zgJZ1SsU477
m9zHWanlXpvCCXACkImAl4SDQQSxXdP/cJT5SJDxaZ2B6o6W1fXmBsPlweCkinjUQ4zXrrD4gDwC
xriNeLYEhfCArdHjFT3iDQ5SKs2KG9yj2S9WBGdwJZxY0o4MmE8VKizMvbF5UaE8FTvMDsNdxTyA
jHDa9MSilXGmTO8rmeUrE4DnN2m8YU+fu4onXo5MgRow+WC3GyOM9olWUdQpgHgswzLJl5Ea3UMy
G2t1s8IiF3pGP9IlyCIYX8xS5Yt6UDEZfEgB9toyLzNhId691o0vPddiGsD1pH6F+hEoflwbBhYC
t7x3zB27sL9CsPFpx/HiFwFppT/rqLioPpcfJmZjwzM/BwOmqTTddynqY5BjgkbIRlTarcIlr77s
ZXVroLgo03e/WqExCQ2DHSqTyHI7YuUE+CwGOtxwtvFmim0j2xLXTOc4u5t4amwgochRYsyMC/mw
Y6eRyo/UbsCSAVOxb2QZv9e6ryRAjxpzWsmmpiqs6jtkMK4az/jCBS/QwDjXeyOkPPn/nltj+vdJ
a8tQnRLyGSdQ/Rll2zMIAdsVj63AxzHfevUdmHO4mXp3EE5pyo5mfyIDnIrzUoKZ6kfFH9fHVQnb
w9tn8thiDygPrklg/S924U+A4WmWgY0JpMXLC8AeAImMSWeblfbJGS8h+t6XlrKtr588aj4nB70H
9A/tznogSmnwHb5PWZZbJEwyXQnQ38W8qoQGdJ3ydXnUh92Z6YPrfgK38i4feJvm2dOQF6RnyZZc
2YfL4BjAiAFc7p/aKmrrDIygOZYE9oYY6ELBzceTAHUd0iXTtbKWbKSqNgrsRv2wDFdiUiLihFZk
6n0+hXsuohV9ccdwsHOfSRDsRJ7HtckT9GTtn6gUl4kUvQH8/drRuWx9993IMivMM3JthtXexmPA
9Fh5C9FGM1NYVokJ+Pf4j5gcweCSktKefYg9HYmqZBpgk7NurZgpjbY4K3TcEBrN4wjiapUEdSK8
TpVLvpCnoqhaZOMahu0OkNJ4IfMjtNweaHhNmoo3cpRiUeRqQUOZboaQJ/oX7W7NQZQaa9vgVUOu
AKdX2jCtIU9EwCJrVVwbZlzchRRarSMaM0JgNK7fJHb2YLDKv4Is+cMd/NtClWzaNT5Xu6e1KSi3
6eoGOwvlSFELsRUAqeyNMLdj1HpV3zZF0+B53SsjpsYU7VjXpJ+aMa5c7AKCNLNfJywRDFVzC3td
SaK4U/SQ/g8+688UNFUJ5Eqbh4/OG00YtCNsS3NOp7dzvesgBHIeGttAms7+zvr8PFOWdGHg/MaG
QyempwAdt55ndjV6s7UPt3Uysr3BSJHgbnglJaImzkM1pIc22iq0NmPCr4yxsj47SzwtgMq4erSL
ndmHpkCyLxLbXx17gx0eTkIHKbXpd0p1cgG/SqzZKn4EMrVzM7mBlsk9fFAeRAL5oqyt3EOWogqY
BT7MLn044RGNSn07EwjE5XX4t4JHPooPoOThmTZEazm0Z8Z4BRm7Pn6G3+5TnQ+bIVphZ1ZDP0uP
+AfFrG/lYL7rD/sn6RGN9oLBjZnFrs4017eZ5yFtdTVmmLhoWNEstiGscCvrt1PcCbuUbN46H7bW
49BAW1h63M7FpmY8loDXvuvwfmbUVfv2D3soHIi8guUl8ipO4ftWZU/+bVONdnttlSb1QfJU+qT3
PLQJgcfIotcew5Ecmxkr2coaXSQrnck+u62GZW1Qf8RHIslzLVEw6/x6ixXBYBWCkdgkKwMs8dxy
GR4BFSQYajUKCV3B4Pnvod1xcjPRLLk035UxEUxQQn3AqHEtiR4KHmbh75CSXoZaYyJgifPKT2x/
xJKBn77e1sL5TIJQhojv3/h12I7705ZB0ifvmBjiYl8znhHSBGtmlNl5mzHZpPxHuf8CgrQClCi6
VWmCd1PU27KkTyPtKmcP4MnZsAvW/VR9Jt5gwSJC3OXBBcqz2H0TORNIsP5bRSzCVfsmqIB38wF8
Za7BJZOkcGv8tZCdCz0d66u3tx+94HGcl5NdDDybOs9xanjc6Idu3DzBCw/lfbV9F1+4Ks1v41FH
FVVDkV9FMUPYv9wG22v2pTB68x+yg/A907ZzTT7LPSsK1baTvJeOXMfXIIKwALfgB+/jNF+29+A4
31/mmDRPTZqH4pICBOyexDdCcBBYzapVJBh6YU0HIFpTl6rlfEYvIVfhRoxQL1zmwsaG+hyyhG/P
KfLmqjjoXuckHNTft5xAsLjxo7SjPwSmEuQmGobhpdQ6xh8NNjyiNBhBlEKKExTkpTmkjKQ8YIg5
0JIpdpllTTnjadyqhcVrmk5vOos2iPOCHGMNHtPntrtknrYuX6nG1OAZKj/f1qda+6A/uHbCXUCm
hzPAdQVfr9rqIyGdzIpJ9TCngtGAL/AHdrE2+Dim/rAIFvhH3KkqbQJMkCPfJdQnP90KHfTWiMTj
d36Fe2tiZ3lgqfgbqS6oLkuC9WKox1UDUojdc+rCED6MQVLDoesm0M3stS5XeJlmFvylkHMxiJ1I
e8nYtArjqmkZe4abvwbPV5wmwHI97YfiWEdukKtlgHrQkcw+Nesz76jqFE0hDvw8opnjwQH6FU31
4/zC7hSvziUnAcbJZVW4egK7k7Lg6+8RMw6lu9XTiO3szSV+HCmwHS0K1fOyzOKSDGe4eeYeYRWU
1gwuMF4sYR1csOsgvP9zh9AkW57gwShqQrjsC4fZvkGEYdEITjKlO2Via+iBrm0iw8Gz7qNI7ayb
awmeOlaYToWxP3kJE4nk1AWp1fWguvAxBxjxEsRtI3Da2nFbAHXGv0imZmyj456I0SKBSILLjWRG
reFz+KVcCGMLESIlJzDSPqfA0Ynf+vQrPZWV+wZ4QOpuxiVPZxs1/5MaS+/YaEQrpXePWurm4Q7e
3kBSs8V4FDtVhUHHps6zrxSl/yOwvxzy0g1YkydzL4ykwEpV9Fgrlz0vvxInWKq5sHW9yarsZDVL
j66CMGBle1JpK82P+58pOI/eYG98grxwBnRqsKu91a6N/snqHUZr072bq5URCkPpFgkGQ9QOm7fD
xLmD1y5wbgiy2D2jY5xYrIO48dFUwTm1oHE/vrmDhfvHnNIBCLk+hjgIF4LrLsKQUw71FvJ+2mq4
aD+qIOfkumX5dOVt932zN7MfOoRCgVubsdp7x/hETTbTbzBoIqjgZ9p7cbkn5bgLXNGQDoh5jT2P
kZJvCWpOXkH19Tbn7UT2kgHRfb9mroxX/cojV7SY47AJMaPB64NpmyJ+HocvEeceCmEddohcTLMU
Z2ORRoDbz7UyaUSerZvXeayZ1sRpCIIEIIEvPzbdTmpbgJYM3qSlL/VmGffpNR9c1XpO9QLw+GKz
94PKRLoIOjf1Cl9ovTOLwfI5BLm9Ykx9bd688FoSp3Y7t7lW8oinnNlfTi5wRQXwr9yWXojRa44N
vh14ovGpuWuENlVjlWcCF5P9p7EYUM5/4ZtuzkUxuYWa53spd6iBnZhMeHropkwcFpeZ8yZ9ilHX
O5d/CGEVk5tc77GDQGBE1/NkyXRBbOPuo8i7Vx0girqA+Rx8A3upybaa675yLy10nsO3EmzjydDd
p3wPJdD2c+SlGKJSvKd7tiqGPTFpwS0uAJTL0xTZvTDs0IBWFLrx6eT4sBlpVQxK8fc50WufbGsJ
enL8D7fDzh1TGV52MJrHdEpccilXxpLo822UcybTrAFlDPy8mcVGkINkg9uUsp1npzELImMwK64F
dK2DjtFuNqLq0dd2WaJbidHrjpJeLh4/xYUFHGq2L8hljVNdauiSx4LxTKivQrZSZrmEqPxGBArQ
3kEWyHPyQttl/RuQx0zd96+s0mJStBX4jze1Aw1Kl9qX9wMyqEc9vbMA6/dXViqZUJkzgEpoh3cU
7CwA/EHdX5RUbRnJptOFgfmW6Q8dwWP9jW0820IB7q/25dbr1ArT4pl5V7UDTnEIPRAg+zZoKW/+
luDfxaoz0T86APiXd7G/i2BuF6aftARL7to+LN+NzXCfeJWl97oeY05tEsV0UkU24/96LbiVWByI
TNtZKexVXIRb8+h/bta/gxS7R3ch245cu3LkRBsQrIyzP2cSFMk+uclyodUGH5ZcUghLwjn1znZQ
kKQzSjsFY5uESSgDyYoQpEwNyoBigN/f2EfzT1oB8rw24PnvYV05G/78slf0DrJ2Hm/i1DGi3MSk
j3POY4umRDLlEBF1eqtxbhN/wDVQSS1nAcXvf/ymcebDQTBFHBufds6TvTAe+6tFhVUnEtBykSFM
F1G3ZSXor4cDK+p2E67eDJ8keBuxMwwx94uA7zshB9URjgLnZ8/uGWmpF3fLg8qhfIpaRiQIDcwr
nfdqHnGny+ejSjHJsz6ElINgdEGp3DxiFOR5pI1lK0625Eq5/Mc9R0kx1ej4E7g93PbQ0vmC5Sty
Inr89eaFNBALKonkr6qXSHJX3BrEnZFAbN94TCxgrqBltPNZjiQZPZELpP0jjpekTCg1adsHQF7s
XWaH9TV//8jzLouwfcdKEw+E49ij2kBiZF3sBm3UvO697qVrmLKR/jo5Mt3+S08/UtgG5iTL8bQp
bBvVJkJOCF2cID8KHKnId1Ldn5MvuM590Io9QqssuZIYz6KgqnJ+DW1qRzL1vtJ1Qn9WWq8ldvfF
iO0rUgCz42HAeSzv1t/he5IZggGGDgi0jRKwXYb3LRBBIput33/IV5iEOA8CdBQIO5FkPK/bIg4v
IR6R6+532fzF4N1jRNEdYdEKGMldmfhNToTxQbr2WGj+UH1woS239l678L9CswyBZC3YCBnt3nfq
BWwssv4CONKbpqzFsGgV/fqIBJ54eb4ik08y2qau7fKgep0S7nZ+5eej1rb/L71zs6t7DVs1TnIH
Ai4/UXWFyN3QrsHJTL1/esVAPepdxiw0mHNkmckr14IIWtoSa1EBueqh1hOUcA20GPqBoow7NJCE
PuM/rNw3Zsqh3hgNKVYLn1etxINdB+WCAEt9zfDCuhHNMuOZi5OkXTo1wymyj09VIDyiZPkFYicZ
tACU7sGch5wHjpHQBfxSGuITezc+t9mm5QYcbS/RTy3/7hBLC8/dPoJkX/rBElFoYb0lpY/lsm5/
gYMfYr7QPEZIkhTY6hKBLxE253NWuvtTlcMQFffxNwKf402D0Ki4fec90I8NuxcVzNHQR2CPrX/u
vVoLxoXwW7bay0DQUGF8Qhma6VSqpDPuE4GYmeCxgzykqW6TeDzg9jVRIwpEQ7EPii0kEeMYaf9a
AlHz/lQ8bp7A4N9gDW8n/YhsYvYIs7i/dJXU9VymSq1h9aLjnvftSlDGWfLe4QxL4kW79xh4+H5j
G4sKNl+EFdn21lruQiG6FBKkaOjJfOvOT01bLpsaS6ocvb9mHjkYfPmcSTULNyQEytV89RcMQWmA
t3mG8JekzIE7jI6m5/iZ3kv8CLlvWtFGtQBXPSmYSJKlWTryeSBf84jLUuoEa+ZVAQub3iK6AE6K
3mJ11LD6gRuP29T79BYTtNZfEIOty6KJxFZy0c76g4eTUUq6f8hofTRvqsAQSYCNyST/awk08E2F
4PDq+JAT51zVq9uNDYfUBbbKbLdh7nzhxeNZxh/paQHT6vw7wEIzMjzFXNMSjDyROAC1MNIvQE4N
VGBcJ1SMBpclPHr4LJ/PfGsemFzbpyj/yNWcAgl60cXP7CsCk4tQ0qBEO2a1OPQFHpjOT+uuFAuK
nUfbWtoeR8/eBkidK94rwdqFEUYgL8DXAxBlun0wSkCQ3eBPqQVq7LBgr002LLenaWdMcK2hMePc
zTZW/a2ttHCOXOJmv+yFNEal1tjl+T0c2HZ6chakhjaDj96k2jYGm/TQzuOSqQhK7C0T0yL7aaoS
uyb3VPVAGbvWzORTp1ToA2eRrBxkAY0B6wdh5afFeT79wkbjiR/X6/Cig9YHNie3kntmtY2C8s1S
DuDZV/UZZtgbEK0OnG9C+BshHR/hXhu3SD3lwAoVDgYUXo3aPzUzJw5mBBkeshHrSo2szHFywWQA
rPj1Nk+RdF4f9lxV7QPhW8jsWKXIAwYYeHGZAobQAF27Z/1zxuBroSZ6hYhdkbRvQftTNo9jvtT5
uiyyE/NfjHF4D+nalBLfz5ABAuuMi/zyJSy+ZvW1Dxg+U50x2+TLq8yuc7/LGunl8dNfGbew9F/t
eh4PQ7O1TA7mQp+ohYMJNrGhhft1O+VS8QWv5kmHImgwQCNJfqE3dSxDoiPnicjO6ahJ0sDzW8Ht
FX3ruL6W2S2KRMBWzrM38kCNWarvzYirsvQPqzUJNfEzYEcfH0dfTJWEUR5/Xc55LanaucjC8hSt
Gw8eEeTHmvEqs1eXJ6f5jASNB0x9kxryZtmYSvniQZusC4dywl+yv7CeV4A8i45s+a1IOD5kdEPX
aG+j44b8+VKfA8P59BUxoKqpMZ8SR65P+GLF4CV0lPp/yOUlYDG20snNSTvEHutZPxl0oEC22woI
8Z7kuvX770fDfQ9NSlwGUj8JQ+tBzGgMbA2g52xAKDcKufjlr8IocNUKoOkvD7jl8YyWUydR+lqz
viocr/wytEreI/z2n+bIg0p7EbyzQvioJNGBdhO/DETug9l2Zdq69DbykKK4VpgjzFrHfy6uop55
hwWbRWl8+YmNWbr/GcYI4Bof8FKlk6BKYQ+0Hl+B7aITGvI2qdnDn6z4F6PGUrWJJl/7fLx08Fcv
LF/6lf+ze0EzudWK17kwuWBZ23WwTSXbrbpgyKY3YOEvAvYBBvpnYobyoaf6IMXI57AmYTHQJWHF
icWlkvoFIOEcsA+nCwE8L4/fMBFfjfMeLYBmSz1fgvmRElQDhFhiAlWifPLO0Hfpj+aXj6+5a21T
6Ggxy8mbmcbHtmT7unab1+U37F/TvGLyzVfPmMBsXEPkcE1k0NuJ67Tt/QnNUjjc8dkEUf8M9siO
EW38+bSJMvaS8+yLhTriVEc3diQP9YDGikMp5dLTnucYepqDqM+XeQcrOQ4Tk3U32WaMz1LoF2ka
80jQ/nN6+p/Rq/gVwTgaBJ9OftfmKcDNQy9xLcyN/F1A7nrHZn/MRSGeITLaXKEieGC2u9hmNlnu
wkowP0H+/T32hIXCFSEHCLVSWRo1QTX/wxWFHL+Hw/xmqkTEtogB83cqN3NInnkQf91BNRIW9iV/
J9XWKXJ2RgTkVmrFhEaCxQeskxQK5GCQVvRUYTpg9t7RPg41jBvq07za16xGAegwjCNtDwbG+Ysp
f3P5bd7GzDSAk9Z7v4M/4coSWVBIDfNzsZe51YXAbbUPVJF4CRJMQZWYVsTQkc52Sxja0sscZSVN
z6829zsR7Nj2OmaB6jsZOlTkJM/vpsrjHh9QCfl2dbCbYRm/m3XM1DWxclrGV+14vUJQ0glFySQM
Wn+co8KOiLcsJ+DHtOp82sIvW7Dkxxy1SBf8a1xvnKYpoW/jSUUg+U44bm/fBJRYpSrjkoKv3rCa
YJxUVhJus8RmhlTqmHDpv6lSx1wObcX1ENP2l0uo74v8qW0Tp5+9Nmzb3tuGTrWpgY/SzVJe14zT
Dp562/265YK8N44svwIRhMJeclpN0poHsLtuHajGvzhRPdeB4LX8xigX6ihGf4LJ00dssKTFpNqG
xY2ItAEqe63fiAV+K9zSIQjRNEP9Z1TKpS60n4bGDLGDXg4B3dv5tqabPSJ/1GY7SkpeHG13+KIF
k2qUmAzS2OW1+B11qnY0cqHHfih/eaVuMSW5gCt35x9oZMXYAWki/Z94MZnLH24YgLYxCjQT3to/
O08uFUWbsIR5i1Mhk/zjQNvQS/5te5T3nFAf78IUBBwOZPlnVbdBIbOPGv33QuElmZgvzaveEHih
4pfgieRY6tGY6lgQ4yVSmjKPp2bPPBcSqb1JlNUSuFFMGbq9X0vZvyA0o24QwsJ5bCivmAuk6bXT
/p20ZNBbOmmBQdkIAKAjya8Zd0kArSYguP2uSNn7bEvGTvXugywCEK3ytLHPSeww2QgaE+1Ylaww
VF6vmyqjYZ7H5Ytgf94MQcNk8Odcv2OaZf+9ledoI7JSIoHxpu5nn0Pcm7at6EIvT4L5zFyo6G/v
3nhcTDqxmTCVmBN1Gjq2QV3Oc+fXkKJRV1em7RZzj1awu5Lh+WTlL0NNqOHMm1BZuHYPN3JHL9c6
mdeh2cOg3N68OJ1qZCgeLDcasV2O3LRjAoKvSyfqtT9VXIomjbOvLJXWWJ0PNhfZ32xxLGUHGXmc
6Wml6o5taFNkjnD8RlLwzKW+DOYllcq67JHB7Ghdz4MpiqtBOs/tP0yidHM/bgb3Z+FXz8wOKaTW
o/uaZhSrsPKEBOHxMpHRi7XKluflPPlWmxjQUHuz9T+vQSw7PVNed4ymRmS9HgacOhXwQAdPTuP/
vC4+rLRloZVorXI0pVOEwtzP60Q8efxJN1MNgtg9UhRYlUEaA4H7ZboOE1sA71rlYzscDo4o68jB
wlQ82FSniB0x1DyJmXoQiioy7wbVQGA8ckLcNCKK5+p1GXhsnp9VfnTKxrpEI4sveYkWfHdmoKlb
aDqZkGLyPelg5QOb9LdDH85R7rFuAf6j36BccQlilC5z8DPGtOXV84CyJvttL78qvrc9NFOjghZ9
4Jzyva6+eORBs/G0+hwVK1xvCwz4gOY1JkG3nJAF8RpI4CAOmkOdbFpDt9suMVG6MN11F7KcCNJY
g0ad3FCY04FntAq4rS4v8bCY/qy0oMNDQvAkC6qaZFE6o85IM39BMDC47uTiUzBLGU3hiXqhLL36
nZHr2QQhj8cMTJazghpP12c3CbZD4dfk+o6YKC5JagY5GHwQWsqw4ARUCIa+dS36brt/vAHH65IW
RIOSWNreiCTPvgm/Gq6PN1HFHptdb6t8TfYnKWwWYsSOiiWuNTwQTU2rs5xH00XPPlKKbm5LranT
qNo+yTTruuHdEu3rC1nLL37LdQ5ub2tEBG6RYBDs6hPUICakrxV39gmRED3zUmpxJNp80rV8Gpzc
mEY80KhzrsYKTHr6ON3poOJGkre1z3fmufrM1Y6Gdd5xH50Uwc2+orIlRIRPVNTt91uLrXGkaiKn
WhiWcXwrZ9osAAQVhH0LM9MbFzODrriVDBNbs2hRbMnhLT3pZcQq21UxIXu/X6SUnw06QBP3rMES
ah/W3DktkAfDn0K4q+sg+hvEguroRkcsPePrRXXnu/7ZTNNXGj12F0pORWsJ4RjBJ7WkVdGLfxKm
Y0dNjjJGofEPuSkGXysjrH2SYG9LkzK9S+pJrCNgUzGckowSMeHeVRWW2eTPceUXmKr3rRgB5JMZ
/iliC8ptVr+63xnKrDtA7iH8OcyBxm2i+5mqoTKob6Si4qGGpawRmfEVq6dqnzk2otAW/njYL4Ue
NOgh9a/NefgU1b/AAug6A4240jBdPAPTwMSm6qCgPl64LH5y5Xy/hb1IwwGZi82Fj6kWu1fQeYwj
OhTJUHNvHEMArfLuG6ofhcYPopBi7fz3pgVZJxLxWMGSD2dMdTfgReZrIwVvRYwf7znuS4zLYrEt
Y3vS69KL522phNCio7UIHq5oB/PpXQGnfDtt4xYDNUBXBIjxO4mQHQs6+k0XUdXxK99rsWwLIre4
Pe3TgDc7uZgYhkzFrRIvZhCZasN3uM8nttB0xI1mN9L/3vypmjAgTW7KztMdBLffed3bPXR4L1vc
kdyJjuOSDa8Tn7G0hmPZN1ulYWymt8u++770fmlBCUg0tFyf5SkkIEJQK2jTKCmfU5RPWPedoq6u
UOJ/wNu9N5pVZc+yrWS5CmodtxkJmlqMcafXl3B0xhkL/yt0Un7wjfgLW9spNJ/5xbcCAoAXnjHF
yqI3RhCx+F8lmbZVGGLYz3Vt0lfbpuOE+yeLAzq7tZ369+a6UWat37hNDyukBkFGqC7D+ysU6sbv
LLh1Ay65+qXDVUTbelhFTjWVwXTjgGWlZo/s2bgb27+AfEkKe7A1ZqChlSUIheNmZgASDSeBNqns
vFzXx5zXx/n+tqch0i6KLKbvYtPFC0iAuWkIUi8bFJz3y0M4UnhJaRNRP6ty143aCMh2tK7YwvLS
H8sEA+PIOaoHVtnLXnnz9qf27hTRtD5MAQZLtQSsSe3yGC2ssSfslX65lBJiaIQ0NoDUe9ijDa99
Q4qh2klraJ8v+8zwW8cwDdfCgvLyhYYeoYcAVN9XQCga1soS7+IJXjSRwtTPVRxIILQNWVFpnsBI
j8BIMbo4LLjl+VBTF9odUep03JS4v4Gc/Y0OpyIzUa3KOTkFPY9w37l6VYFnRJGkED//jwJqH5wt
Am18apqwijyWIsTtVVZrSVLuK0IVnfDvVYoZp0QW/qH2ju/Bp0VJUs2FGqOsXDp6fZRh2ES4hxh2
CzVMKe4EItvqjaSxzxhqJ2agMrUz+uPmRLcrrOMpR6BuafGtngXdZMOJHbxsYFF79cvKNutsCv0c
99vFB+AW7/Uttv52etrVZTufaownJI4p7v1yjE33s5T5KX1agmX1zPptyqwa6Bm5w1zr1RrHJOFY
h7TLgamRh1H+KLi26rzO28rOs0lQ5W360Z9yIyrRgRkQxsJ4e5UJ9AuwRfPcJaop6fq/lNhgKUnZ
M57RVyHhWL9/IHqo5w2WKaRV9r5CcfMUI6RTawzs6TMLGX0HPaQQw33c2gQ2ckMH+34KX6Y6E5g+
CQGy1VTYK2vWVljhcCKCqBPA0x5iakNuJfNSSfvWAJpxERuRYY2bHrKKp7X0HEgbD++lwrpA1o8j
HI+QfhYGsJgBNLZOWK+1BF7aGarnGKSFnT2M9JjKyHvqSWvu+/bmZVk+4owtl3XwN3MhdqbCDyY8
BsxUoAUUHfBleDiGeTLZW5BlLNCUlmMhXsq4kb2TQbXI7qlU1aQ+48KqqeVv+i/0PILOIivyPxRN
Us1qHa8vYCFXi9vXL/p3OIi4FX904+HZI3V6EjsTeXOzGVu/lrJsrjpfvK5lLNHMbrBii6CiqkD+
NiHAyibxYq2RwXISlBSPqMqoiEX+8WWiQIrllbAarCDSISBIGCz/T0sZDhsFQNy6R7/HPqXKUEwR
kFaOBZ5UxXfAYMLu8KNJcdoBmW978E+kH1SxRfRvlw9dkhMMP9CB7dTmCduXd5tW8TyZeMZMBeSp
0vvYWQsJ2KuQNK0wOdutU3TpS7wF01PKYPs0FOIZdRn8Txcr6r9Oo4/jN/HRq1ajdaLzQ+8EDZje
U+eChp35aTmjbSfT5TLSocMqw+M8ui0TdEv6qKYM4myUZ+Tyk7gZFzxvEbUgAsQdUyydJL1X/LtI
t/suOMObb5x9Dg9JM87aw2fjLRD3aehqeYyFHGqxFXFtfUO9k4JQV2kaDq0SbvHbA59J5ytlfMQI
fQDq25oFivCn8hl0PpMbxpysqBScfpCgcpjX3Ga7g16FziNxSewi8ZhybIWW2c+iz+nCumYXRV0P
4vZNavuu2Evgtd6O63548748U5TynsMXx5D5JIcZB0nWLRyjIRzfdKbRAJCloELylrurUV2VmbOJ
aEgRwfuyBpSHwQqJf/WhXFgmw9M94wiUXJ0+JBKQaxqp6865iljO3wpNTFvhJi+ij0w3S37etxZb
iCP95yi9QTbZOlVEaKS8ELixec5CklfUxeM1Z8KMogxU6eZfERFqb7fP/eNak8M18ZAymb45YwUJ
BzG6nhc20d+kYTVWruhLl7PrwF1RrfLeAPwJrizuxiaVBUP4/Llj/5KkVjI1/iPmmHKCKkglAWYB
30RdQJoSMTdU9cxyWbfPfKe3kWna/rzAjgN8KX6Lhkvw5n/QLAiIrIAqp00DeMFG0RZp44rKJgRx
y9Ddl0AQfulHvxKz62+JGSnjeJl63aQVg6/t7WXiV9sEqk49WDnxPuB2LUI+G4QjqrOuSx1H86Ea
DLSqF12LR5EFerxsFq5pH/1GOq6PjgHlLfZxWv1qeQNQMV/QFOPS0dI388TWXakw4XkdJZeYyMbc
CteSfkTIDLU4+8WU+isYTuPr7MFGeKu+SuY+KKg3nZnbCAU+5N6rRzgeq7/IxPcO23Ifcc87J1wj
3WQg4QB+Tzqm2XL48c3/wEB/wjI7QefYkR0gi0VADjzLNL7u+MNKKfzWNwbFy26+4nYEkCjbCQYq
Cu9rUQQdUiXRvlLqqHUByvggYiP9qiHIgN885/QIJgtmQnLN6UrL7HYToo6LE4afBlKESbHuN8IT
NOx5ARZp5TKYtstcvKhZnPpiwBsnc6we/LTooy2wiTuekw8mLFxGxOMVCD8/DEQVE2IFUXFWCZKe
WFD6r2VHN01lca74nuMe3e8a7zx9kmiv1x2ISLbojMLBLz7rgJq9Km+KF/WNeN/xbqxIdcJavpud
SsI+3/QPJ4gG+pOTFXnddUKUdRSr3+R00uIp6vyjWfyvF3qqCrtrrCF7jYFfWuKaIt0sra1OYbwP
YDxUB/JjVijfh0HrsKEtiZRBtJv0iYMMYFcz83bibz9mwsPHP07ShZ/k8N3oD9DU9fMMzHWjFor4
vtAo/+apBIRuOkoUsz8296mfqc+VVmV708Dne0BoZhqMdtRc+jvw7wqTc625qeb+zXVVgwYmjp61
9X0oRVmXvwJVIjkRQY5tDs6PvUtuCtpwYrFZFYfPh7FCLcFDTvmtwRq9DlvFTigq1B/ut8fmGwxk
k77qwlidrRlXuGbJIa3zFDuZx++oluakLouqtHuYvXVy/CjUZouf1UALaDBJvFmMl5uxcyJ5y35d
tFG4DQgt9uNqo5BqPpwOJfy1OcesFfUS/zOpZt1YLuBiQlqIGlQXNIbGC9sidGzyxhKhcD8wrBce
lOre4jIZfgmQ+6nUWYui17dN1ItmppoSl3Bapbe8CH3Hk1TExKPmn1aSoyYTc292Kicz0XjN7QQn
Thv7XSDIYr9hMx1b4rcGA9vj2gVjsPcvf/NaW1YQtTdf3nypssOCszAFan/OMkLAQ6Xjtwy47uMe
WY9qDMGSQ7mOCuqsS3zYQ85DpjVSQSshuMSaOzp/KLhqxJAP//wntHFx+NRJt5p16rzh4njOxdtb
F+XrCyziXVi2bKTVZW9MkWg8JJyxrZm2YYUBR8koj/2CPkRG2HxjOdtEWLVq1ZSRdO8KKICgrehD
6MT2zoSchKRMMvkcLKQM39CgFT/vzN1djaaiRft4bSxWMhwtVPIawA5ZvJJuCZxRXD1F3Oj3yxuc
Le2RdFFS0KziB0SILs3AYkHa1yZ7R+K5VasAj1H60w8BurPUU8IUlAC/71WDrUcXRSCkz/SGrPnx
lzXBlvzDIzXf2OyIrijif9QkVCIqEQceLQ86qtwgFdMEkFftjHVjLa1DAiGBuswt0Q5GMloKGn8M
1J/rK7d3MYejrvwJkR82gquzzVo3PDckQxj8jbggMgOAnx2cW5l+5L1C/B27K9Mq19IU/J6agY4r
FPjU+jSkSxaS/ysacUkTTQ5LOwokvg03VKTlmc1U/sFav0jiONVMTMJRvjkpekkAa6/f+tdGC6Ef
rTyyIDYzm6wsrO/pQ5fn68IO/Ydl8+rXeHmjPWuK+JGiynkj5tYNC6VFlyR1pTiQwTGneZSBMaQv
GtpD7Mrg5cu0L2tKCvgpR28hKwPLm+lc8XmXzcZ2W1VWPL3jkwaNAVLPUpd+fJPQxp9lI3Kgjx1x
cO/cTgNp1cJa2HGUU3pNjQkONmeLBLqQjZ7nOtgtWHhxnh43KTHCq1HAyuzHJzqFuQT1X7VUwK5k
MI8EV2gxeKvYCvfqv+KUtC/eWCZ7Q3VCiftjV2JVq66ogBI48FsMcgu+HSDUbPzNwaC4pOVdbOUN
jRBKaPKoSy0xbrNuxheLtDfn7gsNZ64qhNzmFkA/xNsykibRSNEN4Jjx/beDjVnzG/BQkQqzAYvB
vjwPqnaAbG/s9D7MlnTtcd0Vk5FcCiMxU2XD1bZBaeO7TiPHHvNssyS0BaPZC1AFCmsXwomfpf0m
er6WNvjGUENLpOckK3xWTVwR/hvJgCAW/bUDI2LDu/sP25Rqlg56uNwg5lWmiNOekyHCQVS81+d+
/uYtQxV7G3aqD5NtIlnSKs9OuyqxQT5x/Up2FaL5TguHyl2KiGQa4CU27ib8SM80N3VgUcjB3jD2
PdwMgxNdoF4cfFJt+F58Sfa7IFCUpwwA390H1pwXpXppgz17WSrtUTlfDe+ksBWmBa9F7zt8rjbE
JLPXrLlriqOyhPt/ifSb+jwQR89zOpXx+UbaG7ZTwH0LNjXc9aHZi5uj7QEPH/rNi/zrKQu2M6f6
oCKWrVyX8FAYpGBDC258/UgBSsplCIQoVgbsTrVbrGuotvoRMrl6V1F0pSb1s3pOttj0OBtwXq11
4+ZhwMapFeL5Sm4QkUz7PXcApp681lBIOSen40sW9/e1VYp4Hf34PX/8123+6Wz5QogxozOeyPHw
q+t/zgvDFjLNR6BNZxw421iMuCCTyaPJz6sACqhrXwMpTBamjNu4EhH8VnPJjO/3vl4Y2H6bQpvC
q6vUWSLZzNB2b3lwp7ZR7haesS8M1MDTf1EXHXATBYOcP+rUorRZ/4bJCxnFbh5k8VuzK+1JTqLV
2uMcYAvcvIx+rnJfxFrEPyuHVtQy7PKenonXXW2QM4tLEePwl3csMjVJ9wnNtuyu3PKIIibl78Jk
Zh1PsLZUAa5ESQ2t1sMO1eibi56wOSlSYQz4YcWc3/onFjlDUGI+GlPSRfRC8j8dGtVDSrA7gs28
MoHq51cDs0yLomNalIERL0SRlI31tiVP4lCV94MiZMWIV2vMTwq1Kfpem23JIwyCm09h372FvF7w
jkEYKcQZP252U+AcKYqwjNsXiIcy7cSu9DsaxEf15Wi85BNrc8RPJ4cXWdc1jGoBqMs/090/iL1d
xnioVc35XHqD99sZZerJm4udprxLr+OcmduLm0CEVAV4xCN7r7NKs1nkgZOxwcq/AhyBR/q/UCEC
AabpCCk1Yq6/yQfw5v9IpYqWFDKBDtqsfIzuSTZ7kMi8nP6EF1UAyFZ5bHHG9aNFfusQ1YVyUE7b
t4/dzhiKd4qkHkleggdsbKlHDr1jYQUwOi78svBQuFp4Yo6Lo9rh4t9oCRXG12JdELfjTvbDpfBN
MV5GyotXujJVam+eHMHDcD+mn1rJAjWB8FOzqo4EliNy866nLZf+mqIraoEnd0r2rxBiu7Z42DJL
OT9IgAGkaY1UYSgjo39b182L1geSVX5PWRpbBOi6vH/lZwVIQOy7cV9XsWfDUsYSrPP90G1rSMzV
tCJFFgCVOpqkNYXCLnaELa7IhUYGXOVQJeCakY1PztvGjG+SBH2XVJ1hy7qdIevOJ2oSYTH2o+2z
NQwPCU/c223NmDH98dq2OgFbDfjf+YTkv3WWloAa06EHb7V5oIWljERSFPcjq6+mBkcU7dtVMwKe
z4cJpH+OEfgMzEC5jVi/21pe9SMcacW4/DvET0WCwV4Q3EXn0GiN+pnxHxZAg/umXVRVyaknXntw
2GVxy8dT23R/GabTMd33qvRob/eiWITJu/Q47YTVZE9aSkVgYKh5rRxmzTp59baGZ6oFUEQD4HCS
GVQlBw4XjEfOLGEsRMQZGuyQN9UhwMWQtABg2rFqq0Ic1uHM9F2wnNMQ+b/ioWcGSUs5qraICqmd
52xMg6IYkljchuAD24lXjMekXjOKTrL7GPht9kieDlvxHnEB4m36a49gk8ajf2+7Sl4LZ8kV2h17
AHT82I1hxp3yUHksTihqKtHFXpXkFdu7LdTStlJ5ZC0T3FVO/S1vdvb98+VlGPVZGCHefLLrD7wd
rO3McMwKIeIU6CQDZm2bdr30krtJ+ysnYi+Osc4GV5oULh2PtYGZvEYwi/pn7cnH8Gx2c2z782P0
FpN5upc1M/u5zthZ3M+AInw5XPo3tFrM7ElJKWoWtnvlsf4fUlB0NM6ZMKnKduzvONB5V/5X5Tqy
AT349n2p/f/sKpVvLOP03+BjR/AUCYkbsRwdETbDL/rVx3tQOBtgVrqojb1LZqgmH9ilBfQrOAp9
2U70FsseI6D++5jwxbzAsmuFi5IKUPXDPnEg/RMIEJdt/4ZIjdC/ZDhCmBqd57PLaE6b2D7zODqC
dBgWh6V1LdyP237Alawfqex6XrJU9BhIZFl03lxSPDZAI+0hcfVqowLvCzxZoymJajCjUK2g9ubZ
PoJyh2JfRQsF0bGsadd1fZ+NNZvBga+NhuYN+E/W9D/vEO7tJBVE1In+7sXjXj78uUhW5iTtMQbY
son9I+LhTq8fWdTW/KPbKB3kt1ntLI42+vgq/HWvb/QRPbNmaHD470GfNhautv2HxyAGhApeE33b
Bqt3mvUezJE84dJ0n1vwTz5Yy5F+98BFgEmzz1SzKd3cItzABtZg3taadUAfbapYdxVHxl38GwRa
RAhLd+pxBgaC3OEHhqRqP2V/7fH+CM0rUNks7ML6HmTY6nl/BeHgXxqRbLKGUuOItKj1Bx+RQSXa
DiIzpAKqnhtmrAhq6xU4/OW9WOT+R3A7AkH/89AKyS8F2O4WaiXh4AK63QYux8LY+8ki5c0zQ7fQ
ekM3OA0PeeYvlk9R+t0XI513/bLanrRGWBjwW96noiEMW/yfwtiFkkNhTW9OozsTUGkNnPB1bIeP
ub6GSiXYtc0B0837UkC2ZKJ/rsiBRqEQR1jB22a5JB/puXSdggUYy61JE3jN9BlNIY5TS08wiBNQ
OA6gB6aS42clqW9fzvPfbJxIqfxkqH5/vhud0dwb2ItTxjKHLNzF1makPTFk1O3WUzRGXoKC3vHf
aEOHHEnonCqbyM13F1ahSaj4G+UfHl9c34QJ0p4Zc1vD/eiKGrA/F93IbW5nd/RAt8Nsn8r6wZF+
2bCd13C0n4Ecs/qOdzeWnbgcmMQFdUuWaBkrEBAlO54tj3DO5Vewd3wzO2UQjMe8b4mydbYJRH+u
9aZcNIoTS3gmR0xV4PhheAGFW2wgvnLfPIFW/hkTE23vOfRunKtHUdMqBr3eRWrsxHgCLvkVEq0b
O79c99VekWUhjiSuUL87hMVSsNT/JpwxqZH7iWf0FjAGuhSAi8h28+Vf9amBTcQmu+TKpg+cvfjg
Mlvd7vsffIw5PgJMAvEIyARVMcUl5Xpg20d5sVL0qbke3G1k5fH9CC1oAscTQeKnKpCRNc2izR9/
BfajtmEf9b7OKf+JyxynbqTizswyhk36pwnSl9oQ1xvnTsS/sE20t49mlSV7LZkjehNaj5gbHnUB
GM53U2Ft89H31d0MLmH66vUGEGHI2HKzQ/tMrBOPdlX1+UtgNVvcFUyz5zcMleHVXcgZdKbm30hC
CSJ6qvhLuecQhV6yZFvpfzHDti4Lyt83UR+qhD/Q7CslKeQsoQI9eTJ6s0tF6+eqNQ+hVePdVeSC
gyzGd6zAvqHe7g2Ir74TZisHNO4HZlehvc0xsQVNe0HiY/6LqN0TQ0aoAP5F/pGKKB3Pk85gHFPc
ry/CnJb+wVhQwfG9lWXQDG2lGXl9Hh1xJOWJY7oqetb5Q22QjJKvi0T86UXiVf0OEic2hzx5CoZF
IztT5XhfiSNl8oB6HDU9c4vPP/PPshm6B35QwfG98OSiQqTjnkKsRTzzoyL5yZI2Hv5hfiZWkZtG
oP2qtipYl2xGLeiKy2QP5F4fFPCa1kqdKjLaOZ7MmiT509ilUrcvIYOXl4uZ+MIa0vd+npFaVWhV
2ZM9ghOgIK8hFHr/KW4ZC7/WIWYt2KZ9REYGt6LXhTn8XNEekLfIkyTZDuJPxuXDjsAH5gwjVfC1
MoOAF5DxwMEpGT5/A+jTfGBlxbIWDKidHiMRhKhqpL0ZH9lwmMoJgKXjBt7Crg0+K+p7qiM4zL2c
H7L7gyLNyCW31cnTxkJvX0ynKtJw1q25pygBfu1EYWzMv8TDkcH2TEBQ9J9b2Ehu1lj9aCT+IV5y
I0Nw8FRmEZxjdG1w5yqF0PWJAkXwWgHSd6xq2QEo43xWPx8w5aBYF5nCjBdx8IfD16gWDA1Vq/nX
wl1Y/wKASeX+iUz+BNOd6D/Znw546OPBEyplU8obxANMFrdwuirpMYoOSLreU0sFeNRbe5d6WqBK
wu5H3GfN8W/UVM5kKFDJa37EpxOafvuT7HucO+kuf8Fl6lX1M6HUXbuMuSvH3ypqKCUe92Kez1vk
0TrHUdmeMxnzn0t382LmZAEaSjVKT7tq4h1UbX50ICDB3JA4L8VgGd5cEbgoUwmQp+pyMhlbawec
Eus3KOpZbWd1ubjCszYUEhVX46xZiUrUGFXTv+rhMzB2Afk8mz3rVR0cEDT03kvOxYjPjLPhCE7S
Escd7vYcX+3B5k36KHvaYWyVJCayfeUC5YOmFwDW0Ae026fXoZYjbrfPGJBnqGVbw1tqd2YOj6zx
8gELCwz+vMhTajNuKRbuZ7C99q0pWcLndJkRu9QM2euUD5IRuwNgrBQpHk5XGE1DUS5UjKUevdau
yrhn9A9x6IwEFeaqIOh0aiXKaV6o/PZGtryV9pfyPZ5FuTBkg1q+Zl1Fgi6Dtlc8K2gYvwo7nimX
JcTIZJRz1RaeO4Mezub6etAyI3UixQydYwFqmTUhxsp8RV4gTqposx7hxhpkKWJ1IWDJsEDgEkIc
az8jQfNwdvxtiElxFsQ+0CVxKDiAk1rlYUZCHQmetY/Lzjfm1Vsmb0dULn/nsBe1vf4W/Jtp22zR
ub7alXKDCIWT35DJawibKkkZmlbLjMt0r2OPZNUjObnXKr5tEBqd7E3mQz343KzFiclPqGXnw8gi
13rCMF0a0QgxP6zZLB+Z7Aawl8golXZ2rYcMzR8KupngSwqxwAQBOtvRof+ebzqDDsZhnGJIZ7xP
m+40/HobCeIZT2T5ypvWoyIGmgpdx+q7tqUkGnZyk2Lue8m6gzdVoDTWVb2eo1jc93xX4rVELBKr
aCtCnwOgqCsZFYac2nQqBr9kE5dNEWSUXl9VKFnqo6qf8wKjmPj4iXaNm/2iGITDLS6oetO9YMLr
A8HI9hOEM11ZiqTgKYLlTpRkOfpZ/YUgN+EfWmCIKAdyuJoxa0uKXtjFGRvicRwwg6yCwI62Yt2U
khlzOK3v4Da24gti/9Z9Jcom3SzzJs4hj+qbd5n7MnUb7jmkYovPOGim1IL2MY3NWKJq8gxew+hG
c7clufsz4qOgcr49Y5eP1w4GI6QLiaLr5L4ch2t3/G/YWHlMZFlmS0Fq51y6XS4cd421g48TgtwU
Du0VVMNrXfaotz59lMiJRSnPQcK+YjZb3vvMWPIaw51hzkwlkav9jIbeDsOLsz9nFqiHV8YnHM/o
MLiccJc9ymQ6u3Gp0ackKjC1QPVAQkN6ToP4UmqaX5WtNhJ4EZnLmc3NRtR9MaC62AzQ14xeWl/I
2sVRxbGkoNQJCbb8eMjDeVcudMUpgrItsxDcipzzOycI+vi1wo6Vvjy/08WDk68XWV6XyWypBbRl
hvLO0iP0dllLewTXSjZQ+efiP9148uS5LkznJiNzKJ/sYbXAMzzGxcgfKdmi5hJJcZSBpagA4t+1
2hpPwZjNMXUYlKbhVcWN+VS96EQ77c3Nq++iWG+x3mIIz4R3BvxWEQM6Dkg6E/p6yVjSKICHylAX
lOZopIpzYxbkEajMqAxPJpqQYD44Y2tZJx+lrtvdzSYmy86DQRbXtj6vzTcBigUMoN2eYGK4W7LD
Ep//Q8il68e7wD5fqfIQ5gTWO5lFaR6kzRf99B/PJ4rihCyMJzVT1Tcakkw722gym7GQyfkHjM/Z
4vNISpff6fFSM9SxH0k7cM+iQaqpMhT4q6MMrEKo84ul1G3ZAEe8eE0WCmOuLmYjoxrgTknx4SqZ
Z6CnWwZWCegHklndgNNQHY0nLU5eqaYGCutHOclWabnVUrI7DAMrL1M6QgNU1tbMTF8gZQ20r6IU
tW32UlRX8Pi1LCzW5W8iDN2nNGeAJA2xWrfMzqpomBcCsdbXWpmsIIImu9TwG5vL2MVsboC0to26
8bdki/olGSD9/JV1hzmCePK/XbfCCU47w2mDi4wZVhv7dhDFzGNqfl2lwzuZsyoiH6ov5k7kzaCZ
j2bMhQ4GDbzSFAQjLYWytXgVD6+FMyK/uB18SxVUN+TqYReT6w++8KNuHAeo1nhMuNGCJEdSQoOn
XED6QdU3dwnR35kuSTyzHdHFtvd0zf3adpEBn9/a2pziZ8L5BdAf8c6N5ClIidWrHd5McqQ7sr9C
0+jN7d76oMXIPhqmyNfSC7QLXU605XY6Aq+Me6flQ7wTXEfrgaFQCk7krwIdjv3llhQI1H2f5IMb
oukFLHCYsOBOMKJQJg06U9VaA43Dg0bLJIFh5Hw9hAnRq+DkKsooK+ksQEmEYjKOULdQzk7LVtRP
PTvpQKF8IjHfBzDo+Rn74/ZXJXkDT6e5dLmGpPgHu08yJCw9LuOlTM/KgA+MakJByeLsln3CDz5T
nB9iOgjIdKFWnRgB+bc+9vx1DmmeTSZ2M4fBqfn0b2zc2swrfCwpkvGqf13DuH4ZD4m3k5lgUzqq
PhSOMWkenjZCXWorSGMRtwkgwqQP9hcdDYSXCxY63kbMbrL6ZEMBly1LBAdAkK0QA/Eh330atar8
UAxnLQuMgZMeh8aW8od3lGIYQMFl46Mk2U7NRBysUhJn6LPDaOTsN+RHqpePGFQDk8O50jfKDwBo
oIk6M1J9+2t66XqOUnfw3k01/E0UQkx3qfiA9XfVEriDgTHffsXT6c5dca9RCpbS9+t0JW4PyFmN
yGrHsyaAnwu+QpUhyW/yPGUPWwt5upkPOIPxZz0RJm0lp7zek7g9P8GZuGhDtOmYlpXohGQN6xr8
Xwh2WkD1WOlvxzDecht/1Gx0FEQyiN6KZypz1SL/z8d4L1LsL14TbaZtde9V7xzt+gID9nCDOMOs
7XdEq87MoWxSW9EaR/op2njsd244LrzEVOXeAslSbm+VhmI569xzVC5swEOLzcLr1iNN0zAntFPR
oj/Zv1p5TlpwPzmJRL6CcgZqiJ0/17hxer5Cd8Oudte67rtOKPo9sZ6t0YZk2RcDgdcNW41f+B5I
j4btc1uV1aqgPQtWTjXNr4ztNV49zpDzmU5ZIdUUb+1hkOOw1YBDUOwV+APLhZNxRyPXsJDeg9G6
cMFX9VmzSnQWg+z9WMaKhHdq7Lh5UwxS0IKOY2hXnuxpmmVkD5USe//d85K0VHrHlR2UoizvbnSd
LSsde5uCJ1Xvs7uvUeoImazxtbwDjRyMGJsszXxE0IdoOYJ6w2Jx3j6cFf4ro0hSMvN/uClteiQV
Jlc/sxuXqJdm2S9FPlbi0/NYMRy3rBDJn/DPD58INlzrGAS1VnmngdOZOMn5pNn3nRKiWM4hwkX/
kd9O75/1TZXs4xKB/wfpdVyQsWGp3rG3pI6IXy3BmYK9pjPzhO6vpSUV5QtkQw/sS6IcsjjyADoU
/fqKv9+5D4gFCAf2BCVz0scz6PirP1GpxcrEHUGoKuM55z/XFnP2xmCXtd9EskBg4AVV/vLJ5/Ao
3W97r+6tID5Wa8ryLBgLfR0MzxoFqR1dXHbOlAL/BqqZB2ILPRhZj7FMmWadW2AnE9MX/dt52Tru
oyTgBn5n3JUcjx+xmBlqiJvOPkejQ98YMyU5V1ly89qZHmz1Jwc1xuAimGn7QwsmfVcxhYDtPvYf
bNDJYRXBsd3XD9jouk5i02aLsmX+RyVz0hrTjUuEQSceaZXTvQYFqdM7VYaaDYsFNgeQCDDqB4LH
l4xs3Xirpg4RNoK+vpzuyMf8+1eiy6FDwMVZGeQ+BujbobxF6KKrDqIlVlZv+CpDmDUHbWRnt2ew
SKaxdpimcXIoXaQ1Ps9BsEJEM1a5G90S8A2pMu1e0O543I3rLLDHEP0a5AyRdmJVMCK3tebM/Izb
FqONItBU+ULnk/Jhd7lirwfT1FIHKV/Grbh5IEwX/oisULHviu39rZt92peGRVUuTF3tSyUl+pwk
nu5CCfqM601pcDFWkPOdoq1Z4OJXtIUqvgSzTc3sZoDAy+mY1m2WxiDL6rO+DG3FG/K2xpXSdy0r
SnZGw+fpeflCiCyN3YkbJisP8vjIsIiGdeE5pxjKcoSwEBepSBOHplZzoMPs9PJNg8caVYB3h2aB
ZLJ9ww1RaABP9Mx22729DJFSf/HYwINjCJiMlg87KQ0cyrBkvZtVzQm6LwkcoicATq/iuhEhaZBy
tsOcxq+YYV9ufYge08iS7CXqImOhAoAHb2koGLshYxaz6OlVibIsTpaTtWoF+v5+lzl7572cheh/
cyINSHNQyRwOsVazcluhaHK8WgoEjdruwcwMxoNYe0QQ6Q+9vXJQbnjAZCFWtrK2ADqCw9iiPAEC
SpdwxK092DXPmbkvE/alY9BNnIbsCGiYtGwmGa9qLDTQyY0No3bW9nCP9RgY9+QcgseUQxpm5o54
jr+RTDKhzygcz9O3XUUaYJTetNxszrslAZ+SwimpG2htrvJEjBwBSvfmQBSiFImWa+VqeXOuwiTC
hE8y8Xp/Z7YrNQzFO57XMhWcHloRdwdEXgizygkbttKKjqRqyzZuLlm0rQc2Q15c7SYMaP6OCOhK
mR1GWIkedUvxnjTO9cwjwwaDjDinHpwJkeUnU5cznYxIfZO2aUHEwKXkSx6NBMgSxxekcwRyFCkP
wE2wvfeAquiM7hK6+gF4sthCxBrBur41Ji7nnZKK35Lwntx3usY7Mq5isVy6Kw2RTY78YqT2ReTh
FoqxtYq8nVTAx5byHnQTg8EPNtXi57kKULsgw4uoCyScZJ7lFlF/2o38d1TFnv7AZROo+H0d2vXO
i0Wp32TTSMTUSEMzeAH7WGGk8YDAr7luvdkbpmvFmjPhYbc1lyFvgpefXQ4ZXTao+k8HkvhMfPHz
Pnt5w50N05jZOJ8tfzNiuFjpr/KDSGGJGYzRYSIP4NWgBzfesDtpWwLmR+cxO+qGP60dOg/80Ec4
s/G1UsKgZtlkHuDCEWdJGj1QJdVilqG5GIED4HNg9rn5b8yEuPrswrkYV45N9LCNZoiGGc6/98jN
tFO367ZzTIE13GSAiQpZJhbWbjcfpxEWE4P/mpO8Fvm9utJuE6gCmBm0nag0GZNLqSfI3Tq0ChVj
75LCMdOcagOnp+yFUSg1vJufkVNIM4wcvQ/B7WCdHN2yxXDwtigmlMhwpj4pIfxT3CIWqttLVWGq
qvtyTwOIcL+jkf/Q51uK9UO2Z0R3dx4Ou4ZVaCeI6wRLToubI8pAqze1da1RZb0POs6TEPaFH8ac
zaqUzLv3iyhrVBOaQdft9xpz5rVeonGwF0Jjpt8+ZTZeM6p3voVf7WBjc4LsVwKHel/M98lNhILK
8h7VWgHzL0x2QVpQXt+ti0Ao5AUHcTNntn66a0l0D6rngNsheMxN491Yg91AoLd0fV5+HCT1t34N
j8Tpcghs0XiWwJDBvn4ebAjTjA07Ktilg/QL6g5FP6rnqSmyF3mlWx5oZIwnasQckMvTnKY4gV0a
c4fvw97eO6FGrGeLx9TLd1OVlnrg9hT6Lx3JqfiUqSDt76jVxbXLORwk/VT2eV4lgYA58ElI2d98
Qtf6UREHgN2st7XlPsJf3o2v7YvadPe2j1l17Z9B4PtiXup/N0pegqzxwmdaxmVwp2LH2qiKy8ar
ycfF+fKjVziRrtR2fv4pu2S5iDy76xLJjX3S8s6UeUnIz1KctVLq+N8P0aYKwhHny+akiNBKcwgF
ok22IucNihH4UGPTKuY0H8r0WyqZkkIBmgP/kk3kSnszqRJPFLUnNGXh7BHlnS0QDtmq7euuREH5
EwHuEANrBWxHftRPJMC/YkMzZahb2BVW/V4qZjZ4QaeO0RJ1e2JQ+7adPEkE+4aBIT6IFHHJlu9J
G8eD2mkn+VBCmWnJ8+i8FZjrOl7gAD8tZ/lUj4V0HotmCzYdD8urwT2m5o3TLLuX9Qv3ev0mL9He
2e/7NPI1gvBLGCVbI6IskUKrXh8hyO3jKejkdaDKXTtjLrzRGbx9zcVQpgIdh4QtQqmy8YsOEHKb
rN+LngbT5bFtmJ4lyOe42777/f2mWJYRTrDNACACsxddtDuf8B28eUcYGm/sO6l5Sa2rZv7tRxob
9AZxDuSQAiZyWzwBGqoIiiPEg701cGPuoPDn9/VP6G1FJ40wHf0dnpsW/Em0gLoJULojV44Rb63i
Ay2ea7Qa5xTgTLeL7dl70EM6QVq0wtg23IepYHglIgPRrM3FZLCakglFbH2pSP6APMcUpWd5GJtS
MvQuYwfq/21EiV+mnsf4ndvHj5XMzoZ9Y++1Su9vI7uo5y6Yownowuoe+d5vQrFPDTY9swTwLZX5
KejJFaOuz4JGBvmqveUGyyADSiz1hXi1jmC83JR+AkS3mube3Ui8tn1jzWV1N7DycQBWYddyrL87
B83e0ksQBjC1iX1QiL1oFyBaLwnbR1xTS0jZ8yVYrvWhySnuzraBkkWRWMVwspti47MCuAXgd6Nx
xchFzkPwgGV0tQ2/6XfMesdoVHP9fnQGaBTiG3x+FpAStWlufziV8uQhIZjoqWKTspX0BABY+V/c
+Dq3FgdHUuB9rvqdkQNTOV6L8HrfyZtaMh6oauS+rz8QjDjKy2rW733WxrplLuDpccQabNBMTr7P
E5VyU50lpoqOoNXmKL3GyyyHDbiYLlczn0wDLFLOzmfKWHrmlG3qM3er9WP3/JEbl/ARWanxoiBd
ESHliVdDho7z5XXwB5AnVeUM5FIyBkPkXO8bux2GQAh5WvSwV+8whf3WDcRcevvlQdk1N6dFBfR6
VxmzFLTSDc2X2FSMNE0Yy+mjzKXs7e8tcDXAnHmlHrlxp1I/W+jzWU51Q+gxRPKIvo8r66+BuQr/
I+fZkV8MYDF3rdToHubQ5VpCUO4quwPQ1+UjFS6Og9bfnqLPbU7KEVK/I1AmGMd56d411OEr5xQF
dkA0dPRr7/1dbaXwFN5sn+8vRVKLBnGMGuBmJWMUJohGArblu5uZeyY+fXwG+mkraMO43Ws6QJpa
Uuo/pBfry7PPLBZTrNZkLMN5Ma5RHDoxlTAXJnIA/Z27fDuxho6jfhzPLelBsrKmz21APekOiGVO
8TppxYWn+l6oWmHCMd6WuVvUE8kZWxJmpb9yqXPNxufdcyKJV/FO++mPwNJgmwkQzigW0O/a56+C
WI7ujtHE6GhUJAkHFjxmRI5Df5Fw3eaFSLkaLjiN5SOyQLvKom+ECsqdMPaLrPjZ9WgRo3UeRvEZ
/FTCeylCGy2iR2XtRFxYwTMUeui8/rV+sUeK4vG3Te5cuo5bS8YvUIWLuWIGwnPx0H3aydOogUP5
IswKJyHF/afJrNHGJQ3UN3OAAYVy8Jtk/0Okv9lirEFiRIJyN1sMvmsAc8GEh7O124ZALQ8rCTgb
X2GjxyLkxKfhT4BWM2FsVs7KxO6th+LEZoHtjxK/yjMmS1xwl56FDHMHX/AmL43eFucl44dTTBod
V6wTu1NiV++8m+dehueyzyJJSqz0EBCM07ZTw37fOGENWKB0ZBs3QVONixXuSt94Lq5AahJ2aYjv
RKYbYDBf3WaPlaL7z0HsLgckAKkdVXBZLDG0NUq5gBztkWBg1u51wJU57Fdew14ndovtw7piMna2
OkqSzS6rPn7W7+seEqhv/SMU7rWuF2feEcAhogJ1s3g/scOyHrAv+c4HH7DNUK4QQQiuxpOa7vHz
9qXeUIx3whB4rl8jt8Uhu14MeUzovhLF9pgx0XeGzyK7KbrLVhE/RUPh2io7pBwCUjNGvDJdS3Nu
4cntlETnYERBChv5UmiXIxzVopENrZ8PMM/9v5vZHZYbgeNCtq/2JIcfGjz/aYdfZdyMhCBGc8Bn
0bosv49qokukrJgEw3zZwwgUCwwAg55x1tha4iGL85tv3LMqviWNUkPYfQgAEpVrfScyyziatcUW
1mwWbqMIoYcaduG2DLoRPs0EmzS0rLwpdCc8JqSU47KWhKj/ZUN7bYQF1lZu1Ar4pRxhsGsuPzFB
FFNq+21wnpDg/i+Hy3sSwXkJo8RUU5Yu+eKO0ZFdTBhAObUf7EwMNj9HHFVAe274xRevrYUV4Kkr
/zbt0fI1BpFKvkCO8myDXfEAWmK0jBlU1Weiv47gkbHmWQ1ZLPrOWHGoE6TnoV/1mKnAMoAR2PuW
1MG+2zORRPLAn40oQ8CYuYo7YSLcVnTVh+hCXUuKiGX9KYGW4pdyMpouYqS2Q+GBPCHAt4wYyCT6
eaa8qCYR1koTlw97kpot+kJOs4kyL1gBWC6ivXytq/jeU4kjKOK8PA3kJd8GMfDkzO0487FFmiZL
7ijgPpn6qUpA9RFbjaJtkCxpXk4pNAhki0HttNWG/MjJzI+c/MpP0u7wlYfnB2JGUJJsG06+G245
hKgoS42GblvT7HXJjzWD/Yvx6OHsjC77EXiZB9PK8beBuSNfL/MahuOKKhgI03oXvRy3CtliRqv2
m5bBajrh3oxNr14+Mf5WF24hqkaZWfjhwI8WRYcsGNO9684ibTAkdz6VrMST5K4a+popkwVxYa+Q
JrlNAJgmP1JOYVb6bVV/JbnIucdXJR6rnGJ0etDDlI3uAfrsjG4fR8bl9Tmc/XlwsXnVWMAEJSqS
kXjkGiUNtffKYtj+gej0fpOoQOY2fhB7bDLB6lMPJlWw0IAc0J5LjRO5P5lfvXLvpiKHvYan/FRc
NBLBpSWhNu4uiaRPCP6Ohq4WLinLBOSDZhSSYCvhJrWX8AML/RKuaCooq+ThdckMRRpYkJK7Dsti
rBtORrFMl5F7hW5ThYyBKc4j54a42bIEBjCYbKGM325dNBYFx0SYlVd9a0jXCadrrNMxI+3oYzJb
tgVxuWSrzRu+T7hHA0H+uuTMOyp/GXtY8F4BcSVIa8B2JlhHz135Wq+kX0thDnjrx0hNjBzfFDoz
OA4GSeL15qKItQPuTqCliZJyma2SVhXuAAhjvV2AYf7q22UquOv2GpmCLtJ5XxHI67dGc4zvVdC9
w7JV4uwcQvOf2vnWu60HGhpd4bhCICXWKmRZuz0YbHpiZNH8DwXsAVd+jwKjbqL3FQy2qJedBI6Q
WyOdOyqb8We2v3rezyvgTctwmuEgucBMFtVUl/L01vbrUnz1J458hoLD5S4eprj0d4XIiCbkb+xP
4V6AfnxldqqwT32NI094O5aRSVlrh1IYTQiRAJ0FwyKV1P0RPGhWUgg6jUzjzf1cOoJ+KFfVVQIP
zwXo7fHeSc5NjJyuPCqUAlLsGFaDqRVFYYKq/ssJu1qHRZoiHz/Mj6CTO9LbZgyA3jwqob6WtI2q
sGryuSCeGAjs3sJ2kwYPmCFOgTGWPCz70EB/xsZQ0Ku8F+xD2cSYxOIbA8piVeX388q8MIAj4lwf
wEhb470xYBoO5DYjz0zpcAOxdEZmGvm0rEqSylLR5XMgANI+GkSrZKgmVSk+qR4dnWPLfS7f4jZR
96nYVZz/ckmMb3Fs+5OdWw/orhW7JTwLK1aT9UmWHBtP6fh6tv/daefEoulwjH19pE5CvolWPSw3
YWNEyEhkA2Cn2h6a28tkMEDZCUAQ+xaPU0lY8JXvtysb1oGd+cV1vlsQmkYTzXMXTwrwBegk75bJ
Qgk4U4Hb5Sj0l6oJ4iOWxOLimTsTj0xRDA3XA2LGkkAnDf6AOkFGkVca9v+DxJfb+konj5qauu5b
X4anaPV6abSuN187N9d/9BlLFAIk0N1023XdsIXxsrrzwiOGqQLX8s1HAN+Jb5RdhyWgncqVRKyo
pKXRac4O9vqAARF4bd9aJCHojw1blEIe/2W4Z2uCPK/kJ/2pAv9hdnNjQCj4qYShlrXEAZUKv2Gz
wV43zv/W6mzRBXYHeNV5MVPXDUHlMmxzoL9PbflHtlHyLw8Oe+7uyuxk3M50Z8V+RBif869WZSXI
N6ej7CKlL7EKVCm4rHrZAlLvJeV6bZfr4BRYBbH2THeiE/qcmV/eJDa2OCBtmbq/VTrgZtq5DMkQ
Kc+wgQrekAzOe0pHkT6QBjyzEzjuyJVuKvoafn+x37wVLMKCBgaht7+SU2xeWiJhMcE1RWndhbfl
0RVvgjtBL4GmktR5b0rgBXSCMntViRkOOyM8AF3YIbqTmE6DIH/dndhQjgV6YQ3yVUn8UEXdKm+R
gv65lwW/cxQaGw6SQo+uFt9bhuPQgwEsdLqsU7IkrweuNAAU/IId4CHdAUtHifDn4FaQ1R22cbHj
0I7EL/MUXEErzIXTGrnYBoiQgVHqsFq/ueAy+Y17b/z0rKFYPR901wUxM1FjAuG28IrwDkMxCd+H
W6fcqbMhrIiin8fWNJ6273G/2GVbKKWCgqn635gY4y06C03dWWZNpPAyqrNtNO+LwLOIEZEZd08I
LMuX6udWCvhE2uv4DGvFb/qioOmwvx0YRLUYN8kXEjXk8f1aqaLPS8NQhhbMOtTlt/TfJ5Nw7lCt
34RfbbI3EHc4GjtVQqe+VY2KPkcNOifHD0ftSO4q0s2067VS+KaMtD5hnEcLEZOv/D5BK2/e3Gg5
QZ0nGf0Mg15UB3QHG9IpyC6ldNcy2b9swxAIu1Ou2mhFIRGLxoyjzCSCzBuS/6+hPiJ6gdVBMbIL
NMuWvaLu3OCun46Vo9D0UbzjIrjzMmDEKKQk/dOD7FwycfZR/RWlgdR2+l56csQtfdmXxX05yPu5
EReP78HZxCUSXYe36wi1JUH719QCvQ8/ogOUvKE4OA3qYLBO7TzKSDmpkn7n2fkgCKyGeHeNho3y
Ty4Wv6mJtGkgkjEJEKzPQ+IIYsjafiT+QGc+uA7GkRi2pcsLhR593shRBGxOzMd7kPSfm9Cflgh2
IXI0AqDy0cDq260vlAiqcrxgMQuorYq2ztProKbNVw7CLvRLAUCTWUhfcLTzNOEqHpYDNhjhde4a
5kYaS3/0tn8PQBYyqj/MxYCtqMaYbL3yk4bND2iASCQfvwDI0JuN7TlTc7d6tF/mA+dX/kK2CsJ9
5j9+JzV4PsCNen9A7dTJYjg0auVDLjnXvTqeAhUvThh4iCOSFKzFRsSqzXvkQAzFQURW4cBGSjV/
wW/MAw/mkaVZihMmSXta5gSaQZqkfb2vCDXPGbEfYsUulP7IyniPocio2s+JB7mY+CUi6sRZm74j
RDY7q4T1LK7nCUvcVSU25hx4jlQOqO+AiAnFn39wF7VCQaBdNFxQuT02p8JO/puUdy70wDfoqTsp
sH49nCHOCyWTCyzyzGKa/wLzSFnBuZnAy1JE1+eaFJRlvH7BQysBNYnbv5eoUfi0ivUoEUg6iq0w
G3NYE0VQjLZZqF7CB0G6KUfs9UtCKV3u12FULzte2BqMfLsbOUR5yMnL1pfWalgY8mroeB5pzDjo
TOg3yBC5XlefFWKoQ4yrxiE5kMpfBIqcimJei/MOGEYtljOsr1EaydErCVgHBFW7tyEaxZC/T2CJ
NZ2XDEAaP1OuR1z2zRZnAwlFvLdBgiGrcZxL7gQvS7b1fXUlEOAzM4ezkZBZERAjWGGdoWoI1Fet
93Jl4KBBN6tFZpCYQ1typ4MlOV4PkUW8hlMMAkoYD8kGwyakLAV6PJIIn+DTlla20teHIomaPpRY
uRu8D3UD84Zv0YWRu7emXTC+i2N9R+QWgLSV5wtBYZGgiCWC9LQafIIPlv7hixHlKsXdQIUHVSTN
jswi1F1B9mRmdLyxnd5grNKemC0+qbTL8PQqaGiBDA4ZIMguKLCh/IVywp3uaRB7arUzHK3wEB7g
At65RN1WcemWwwk6pBrPnadGUfeDXR/TwDtlD+m9CNbqzCZvnfRdKlBIM7WFYVDL6zaupXRLuyRb
BQjGq2uy2m6i7/tckIqCidHuRJ94yAWuRQVVl7tuaGl66mBBJLFoYSCXQFStyMsDIi2zNq1sb/qC
gouCljGtMNJNJcgF316SSP0usCeJ2o1EaC9N/wz1kH34PVfiYgrTgKM4vlK2GmswCDjY4gqktPUv
eGF/PXDFjp1oNMPwYwpLyEnVlfWZKsxPcMSkkUSgcMGPb/xHQagKI3DsGnC+ytQkaF9owPPuSAqZ
yZL2CtF1m0oISvJlODaXIGGBznqIxawHmqMGXkHXXiUpWo0r/oZSXDxvhnTk54JdQ0e44W1JuYpw
rtt15Pe5Fw8UvgAKiIREzgRt4cTghjdAIUM7Sl2r30T9TPBjDSCJrV2rYQiAzGhrC6X85bSifkfk
azHBRKOvHeLdRlO4GsMbdvtzPihtKbmGTMvyHYNr7+8safJEIKXitCwPn8NWzJRfzIfmV3jdvJaA
yKHLXQYc3OJEd0SVnWe0/PioG0jRJe1K1PMYMbMe4zgoW98l+319PL5y6cTetc3xblLOMWLLP80z
u+lL7oSpexRzWNJsxprNIW9cs7OTPEctlcYy3d84KVin+DZmaYLy+TBy1vouYrWhX7uk3HL6stkA
RlkjUy4b9WORS/W/sP8BBBOdfwffTJ57tNGNsRj12pcGeED3J7slUuxk34WBGzln9Y3b84dYuLsG
Q3T4jF9GbqeY3NJIt7h9hhU9rNLOrGi7c9R8etlReegA0OuMl6vlBBVh/GmNAFkER8WCPKBGze0+
kS6cd6O9Cr0lNOKD8PjBwMQ9BD+gKQXfxBLRmXBJmOx1CEUhk7EkM/08b1HLVol2ML0tnLCuzc0l
y2VxSxp4tlPTZwJJVFN9V+yZ6XB5qtZ3ZDeBRdlfVp3BhrO4H2HQZ3D0Xdy3fEp97RxcuFvEyKB6
VtWE1UPNPBkDI2p+kGxwnG1OVAuRmXNTHotN2g/eSUGSWzBfarFogmFC/H+sovsaNTzRTavFSWvl
BVifjh6/iRS359HyVPkKfqsVJ20zkoRvo8YgmUZuReuTmP0+ZPsc6Cx+C0uqx5ylfoXZorWx438p
c+2MvhwbRLKoj/yh5CUucakUyn4tXqBR1lVLzB/PLQAT4muY3mQIoACXPeAsbAZcV2EVVw3JOkdm
hoB6Lsixfy3jEN31BXOmGxqSijUpA7HI04Nj5fe7tTy8TOKOhAItXfldzRATW6CBmniGBM14dr42
fihOKS04+6SwzrtHpwNjRJ2BC9woaAkk0PBONWDe3OBzAC9ewMfDs+LOHFq5KYxJaVBh7DAF98g7
eGX5LTedkoiueIPQi77irqOx0NqadRDqvFsVhDi4LTKEap+kTbqFP4BbwNQ0lIsdmrRndKnN/hmM
lZP6aaIIVApXw5XGdWPpswJpFPfToj2Haw5LqS0RZP3ebXDJpPQHMhKu6BD0DwjHzV16vUkJjilW
hqbiNqKSos2AD8dBbQF83VM3anmo/FbcDZozeZDv21qRqf4sZd4tzRkNmVQRyUZal6k1DzSp0Ztt
6ubdzHRO4sNK6ILaCDn2T08nsS7hVJhiqm/MUWZMKje1BqoRThdiPakugTGNAjVurQ69pQ5KM7Rv
PxRaEfGlFsngK5RHlv3sJHxbsPSNwoDbmb9IFcjccH77tF4SzWLwcLvl00JvdluRYEb3ThoAdpBl
+zXU7aCdaJcC+/fBmuwcreaPVWinIBq+ANJSzwGWlzr45cZiV8rHTErOTwFHJgmE0dTFNt6Fq52Z
onwtnLY2oEXCEzkRtVVRmCgHTcjqytrkhqTJsIHjtCnje9eWB2FAcGeEEjOldHE0TLHsWPsftlZd
zYUhD3rn9UCMOiANHGEnMJntK1o7qbH/y0fQ5WmN4GVn01rOUokoN1/02oMypMre2xcRVC1Qo1H+
tEg57B492apzaIzNHguo63W3dyGy95nG+qtPAFamJ31rIu7+irVqHbtAS4oc1OkRa1IaxDso67uh
AXvGj0b7M8fHV0FMEO8xRDH7AZQyu1EDrWxutjoZLJW/Q0cmCnWrbPfRnoPZD6HX1NpZ9t+PkEaQ
wxAtAqN4gROjiZBjFkmdDidpzY2JGVzXsMzlXZtrbZiG1Z/wCERux5ZfWytvSJ8b6mFh9cmvaJiy
zlfWSmSEMkT0AmbRjsqaSOJCHp47/l3Eu+lK+QhdOfCjpIJSYrfC6HNRG0WUhJkIBC7XxuYm3sh8
WjmyfD6zCCrLxyKwglRXYC+A0nZGI7SwwehsWE/ohKqiahnKftztv09Ve/S6nkZVP7pki2XpUIbl
CUzd5KFo+Ear9iC10NM7+HHbEEUIETr1743VdPpaStbeV675yWEM+gHghjscOWvEQsuXc4tM1VgO
WueTHLlzoIsNO97uB0JB1TVy3yP0ddD2bj9wJKdymC1PRUuUd/thD5kJt2yDVohzS1UCmwuPvqOU
BJFgeNpNChqRPVe6y3aNatWQEaoX256USOTXcrWkaqukUS7NRr9WMmP5Of8NuHM+gtp70fioYtR/
Gh8Qo8DEwCJnuz89wgi4fJtOsjx+dnfDhLtNVKxhT0huRtIO3dIiLgalmz4i2QSOC1Ax76lOo8W/
wlYUFG6wkfg4LereE7lZE/1wyxxyQMYayaVIMy23A5tTS5u3SixDrCeSzhEL2n0Anaj2FewTTE2t
s3Vhwq4K9WirnVPT/EI/tvnAu/n4yG8fcuvUy/BylEIdfoA7evxs7Tz+gQLJIiATFaS07TeNPTW7
fk6inhZbx9PZEeevMW+J0K2q05YUr/CHPP7WAemFklkZ/I/JgeYzENz+vP7iYIncP6ivMFBXr/qC
Y/vaCEuNOft4eZtaQvDdL9bjCv8coEKKdEy22ojPZW3Ww95gfcL9ttIkNauS7uSoaOHKq6wxO1m5
1fveWa8/ItH1Qcdzp6TDQ5kM2Ycox9Wpm2k2w6w4sWBeCxLCumNAC911EthyLQ+robeiLsMW8UJ3
KZW6rMyg8J30lY3xsgWPp5KoON+gyS4qu3DT/Q0W0abWKvOPP7ieBBNQaLNLruGSG2MDASg0DzM0
Sin2BKtnR7wOOTt+WCrztDDdzsyx+DBqeW8AzEF2Oei5tpRPI2MQ/4WBuaRa5Nwpr967s3rFPWT7
jYC0CPr7RyXAEag5WBMr3WahN4sgquJOcksxJmTku3EDt2QcC34eNhupAwicWT9CF25KW3bRGWKk
Mizu1GU9kLtGpW/i0vEbmvYoEN21gATio9s8vxUNSTHCOBr8QXZARMwfC2ydjp7rR/gagKSoEqsZ
9Qd62/6S7mV2HPfxNU9cNfNEwmhts9uG3EgLV4G+JPdWx7m8YAqJhr7PcrTC4jmF1k/X0OGwnKrj
YR4TDm8Aya6qdDLwlQaOTGlvt/OufkDcDrsT2fSrSX3uNeEXht8IAyfxFASca+IHSC+HOvUDWSVg
9DghGcNdClZyBeQ1PhVdGehD+CDYiERATo2HNyTwC5KaxASugRSTR0v8XRwXK/i5Z1IchMRdOcXS
xP1vZFZ/KYhoDx3BGqW8+B56ibpKuUe7vDbtDgiHrAQKOfl5fsZ/MKDd0DWqKXSaopH8bFpFVkcI
TOfRY+o/pnWgue1rzRCddomhtejZpHlTXxQ/d7BbvOLfvhZqxK7NbknfL0/PvVFaUTttgS5AuQaV
VNxbx3ar7yTRF8JjYk/d6RPHyYol3FUTKBB8v0E3/Wh+wKCDTWVJiDhXxFqwjfqIRgs5Vi+nQdP+
NT4T/y0Z0dBT9yY2TV9eL9FHs4HeF3RXwvfXOT44K/HCZlM3AJOH2UPKjiHe5z66dP7pIoDu3rAt
Jk/oHO/TLN+yYm7j45MFnj/BsnN7659dBUEyXfkUg1vCJ5noZO1X3paol6R77ryXugRPH3b/HI3l
uw2ExrTKfHCTQuXtO97U8eaC9Q/+MTmJh9VoPOGXnnPBGG9z0FLevYNgAvbfYwgl3PzPR/K0IsiI
/8U5RXjGVpPcf13ks6XTQul8oVpBH5riyUIRqZAx3v56uyJItNVJbgaLPW3GTjB3IEw2C3sSkZt4
Ng8RnEH6NLJn8mwNJ0Q88XKtomr79l62ZIesVWTaP6Il7FCxmqcOtZmNGheTYbzxwnnMFEJ8DpGC
CgxJO4e7ga0TUq9Mk7vN8xQY9SaRcA308Yj2JBXkCLMvyB0rOg0JYhBR9c2b7ZvkKWGAh4uPZXgB
KkdGGbYzLQZtWBgmpXgBIoDuAxxfgVlgCgwApZShZJlItpvpHa9UElDdpZvfg3c5LQoxLdGWB+pG
d/X3F2sN1kLZAszpDUnf1VvGCFgiMaS8cwaJ8PkNBEAph2aSNcZ3vp8aHkgdonFJbEj3lyz7URrV
KynmVFLfu6Fhsum5NhRDhZmbSKotChAgMHO6Vc1m5E1YdPXDM3hpb7LZ2TTrkgv/lrx6bT242zDS
2PsMjXkWBBoRLBZbE6RQOoZJ6jXsmj0JMqeNze4lB2Wp9EsaigfPv1kC1QYNF6ZCGmZVJdnSaIVd
Y5KldFcxmFosZRsR00UU9v+oaqHiLTQz5ucNx+sTWTbiKJBJwfPduReXIexr1c5VdfHk+gTcWyl+
0y2gK7GTZo+qLR1j1b0iu8I0C4Fr7gBNRiYCaQuJTiH4egIsQ/Ml9zP+1yF8Bk7K8FuWjjHmH/98
m7fE1j4o2TAtvRzZhF3CQus4deKHN+KuDLC05HXRE/YfeY9r1DyUAOutRXOCqBGG25fh/zMm1dfg
E9IuktLGuDc2R9W7OA7Tm89EgE7YD62T35eUP+THvqW/o+RQlrhbZwcQ4jFH1+lRl2XiDYwxJw0W
ejFdj53Gwaj4/JW110YqFnQcReFS1Zj5Vtkh9QA5hTUyfx9hLsnS55tLKdMEi3ystplxv6CofcmA
iVyi5/WvFIaaywIs2HwgB8DtBl/r/h3j8QoCpUKoMPuaO3w8yvJG5TQyuyhILUUzSUOF2gVio1Hz
Q2Ks1tUfRdP2NVqA9/VDpn2RmpLsoArfItrvmdTpvndyqQnGqZX3eQHvLh6bGuy9oUtwl9S37Bnf
Zb/uZGjMkiu4/rbiO9RAPzqHG6naDBs6399PIS1BdPOo4cE7+qEc1cNq+zZgPqq8HPhA5Q/Ax94w
CdX2CooZrCsBBXDAb6eFddv4O8mHZ/irX9dKBGbH7pvufec4hRjPrXeivhMn6SC/dIoDru8pMiww
0mCpxyrjGz3YN4CMQeFdUJ55h7GA27LWwAGv0onPPdGrh0a8swJmnimZjngHUuTTfjRxCQJiImMp
hHAn22hbSdmDHc01doqHVDTXCTM04ynnefRSLEDwb1wv9F2t8Q4ity59hqApDGUqrqse9bVDHt+H
4YJqrRId8NNM/pTcRqfUH1N12CDSpyM4GFjkRIbpUngiSGqEsWvIkSS1xwlxWKS9U6HPKkxh1BBU
/BSUVioOZ1fJXqGeYpObBv38+OA2HScSd1tC+A67lKThxCyQzQsKZA82N9gGtdOrQjD+mqzhU0qk
ByLpm7wrGn3dqkyvqX4yC+u8G+qGq2R0dmlNS6dsooqPaitE48yDixcgzuIk4fkmv/63UOh2euVw
k1wT2x8oiSxDS0ygSP4BxJpGdhNUQxXzo9GaJD/zbHMnhkIo0+32yb7KddfTact0OK6VrQiEg8jk
ncpnPYwdBgu6aenHw+BLOAImfEK3UTIDpDAGy+IrAJWEAnWmdm6I0G9Bd5VOyY7MxPb4IIDkv4rQ
wAk17jZ3o48PZ9CgWGdiHMJySdD67lJPPwlR0uAHOzwpix+6O3gT0O4hgqlYOu8OHaCbH9MgP+f9
csiEvqFfRuld8IYypvihxvyTIQhrqr54ZWBoHpqH2iWC3qJclSF+y1BzoC84GVbHGTh0kYMaH/Kv
S0fvnlCyHGAVYH7xhRgIWUnWnYu3D40mYiyHx0rU77+Q8QVZDI+Qw8LpS8qMYbtflbvpzDZ4lCG+
TwKEYpdD4Ahq+9i/KFbWEYsf7ZBqwhRf53skHXD2nC8OhucdqfHirSXzfUxkm03nTGuD7DCoVYg9
8Yd1xF/184RCMB/y3zGx3cfp2iDyYVehPYrdEknfL8CZnXJmm4NTXEwuOHaxSDUcg7Qzj4llGFuy
cPB5jrel8cSshnLp9wF9OOh8xA1C30Yc706G7XINyiRJj5MklHSPMQJRE7Cqpd5EIJ1dbtqwTLhM
bX40urDfmYTmRQDvyBZNcKUrJXyIV733c/DQ3EISAqcjzlzD3MT6wOOrd+atUmoa04gtfLETeBoD
FAs16FZeKgE3zriAy9M4LePx3e1rNIuvKM9/sOVax6CBef6skgNH6/OV+hlsfFfNWoXbm+NBAEZG
eBoK9TF1uDPs2YA9JJ6YLxrCB9TVvQ3uiCve57vX2jfjA4Jr3R51SIyd10wXALRPGlBse3L1PV94
TRT3XOVbf7QXdFaIMPQ7kB19LKH0IfrxLjbuTQIXtYqdGHN5oC3faSpr4ayTT+NKPZkpPN6wPi6X
MTusQJnbEmGX4bB+8COnEyQz4AvdhThvMSAjTFJtsbWrZggb7lpWrJmQrkZmjnSwKCBd5kFKkMNF
qSvxHIgyzruyBUFGGmXnF+HQShB+fzhOlMKlxXE2/b87Yy+OLQn+jh+p1gpW7H6hy4SJ/31d2No2
ipsEIAHWVlGwPc5mR8LnA50mP4LrGcInpOe/kOdo5zP3gf+FsZ5Wza9PAE1tJdnzbL1RGmbkWwBx
Rj0S+CgPeUtUpgk7sqUPqC3BgV8m79C3VFWeqjQ5oc2NWyjhVP13VBN4exCd4Q0pPU4Ad+GfWnp/
1dRBdQsO3pNbmUdIaOti+6a9dREDbdx2hFLRCwgLMmn5nUSOY9Mxn85mYCOF6YpCYfAJh8rwW8PM
huFPPXbP0hyrRSTs+K/fo/r7QmQiF3O8LBdI/AoDLpbeQtB8/yX1HvSGsJL54oV7qOSrKtHwezja
Lp7T0opZgf3nA/MetLvW+eEfzZ0corl2emhgi+WEiWnWfkcBnrmj3eAldwB+XIRzghXnUUYpKEiD
ixo/w4nbzZYa0uIrXclWC83aKxWsqOkobdOVSPkbVw2VXbUmHEXWQcgBNB3sM/fBWep9MbO9aRFe
HS1DtHTf3hdaN7f5hqdhFrhogVlgJZFa0MMhxL2ZiDQV0FA/9s2V1PyxFQtNTxRYuwC9yv/0HcGq
zO3BPxVlH5eaXqRk6rO9x9csUrfHegyuiPVaJhNXZAJ0nMKVqxdxpIQH5QDU+KSfQbfhKKoZgmZ7
ODroQzWHcP+vzVQ770obmxqz9EC5HsikRP0+5+5Keiwrw7Nq7NcjdVugRtkWAqmQnnWAZR0cogNN
WdeWmukN9ZhySIgDKZWxFJ1qj6E1D163u0C9jFGzHcuoiXNwhYW91ZLrmFQFP2szjv3JPIPo41Cv
BZR/FCoM+STEK8T8idiWxUsa39VJX+I0Ar/yLn5BUJXEAF/RM0MLu6I3aMS/qYYdrQk9roRM+izK
TT87ogmXNcURhJGKSrFpgfkxXeXmX1oC/kpZG2wKq8Sl5kxCc5fXApsw4Wxr0v/ejV9eLrrluryi
Oh2G/Mr/czQArGc0ViUDO0N2Da3vw+EAoQN6ek7UJqvha+FxU6X8yM0gr7Vn+8/pF/Pnmy7QDYLs
S5ql9s+i+SjPhhza6JW/t3a8C1bBcX1ag3FWOmCtfZ1HKdGH74o5K9z6aER+7vAxR/RGyob6639J
j7qZsAidUqKsN/i/KTfcqn5k2Ry7e5bQTrupCO5EZX/O6JQo9ck0EyDJA3KaTUOCBZYrgQw69FII
q+km58aLTl/txyM4URQefGcqJqB7yRcV+JiU1TXL9/RvZhWBNT01o9dA+waxPNg3kpk6+SbXT6bQ
fLkH1WMkchhPmF9ibG0ipbD99QPTSR3772/S3M4fPTanr0pFJPzksxPDmP1DeEhQupbZY5C7UnLC
lK/zhNOXmOTCZNdZrJVeI10ehYaO+WdsHV1FlholIfmS7Z+sLE33NPCtBBfoeAsF7AjqtndIKtas
Z8tAkeIwC0wNAfjXa8YKS1iHxjoHnbd19f+0SN39/jgQ1wdxtDFDXCTFvmxPI7mY9hPJ+gMqL1cb
NYC0HNJik8DarwqKUmjV+yKS3OP8k9UDUIBs5TXQXq2hZ6W3hjWJS16bvs3ASk1T1hDBjWrQ/kGk
LI5fMDABoh8SqElBx0HbMPDx12K7+e/vwcSM3roSb8GdaH7lAsdwoO4lPGA1ueoNmXlY2rcIXABh
+a87C0G8VFwR9DaoqBup6FrHilXen4BMTVQR7H/ZZe8afEUBZ4kC31b+TH3MCMNZkeZaZzXn7Ybp
q6bnt+FoFIerZu/lcFE/iEVsBkjXTQiQ6gGcZfyTkt/SCz3pkPhQcKTYkTtK26J0hBCVlAVImLY3
NjowgFWSOmv1yVavVByDXD7vQuljhbfx5TZchFa32MIUzKHypNPEJZAW1pnLxbidXCdVeeY1L6NR
6vbTu9CIV6la0wpJczHO+HbmleOC0cpcWybmi+qiaViXG+29sN+pO3yn3UDvP+cg/A3yY54zCls5
2DaVlZHbBDewHX4LbX8oC3yL0FENOfNoQoS9x7EbFjEVbMoQ7JhZZiZWpTq0YUMGOjtNOG2WqpBz
vEbzd2Bej8oL/KEQxjAGLWTTVTNX45XjPmFdDdHD4L0IEleM1UJ5VLBwbWa3Rm2U7INJqoQINTVM
4LHUu9itvsVLcBDt4wD6Yyx/ajrQbwCcxMYbzrP8YWmqnE6OqaHGrRFAZYYbFj+6Ze513F/1lIWL
GKLbkoq/lDjYgFk2E4qGInJNIbBeDd3nfXVil3xYMxzFKTz4NB8TC05vq1LNHrkQZKwAJkiqpAUl
hJX9aj3BxXD6uN+82fK39oMT6k3OIbb2HitEc4IOyFyHc4GeCch4lbyA+SGJWVmtad6AJJF4tCU+
KSlsnYEPC8WDcf0BuHwhTCNtu1vhMC2GPNM48YGQo8FNsPYdPanGfelBTBl8eIHdMrGhfzYMHBCa
mtpd0eUfWfhAbffugt+dELsIcr/u1ngNN+uWCGJnkCRtI5AWzEeV12uyuvWwDuIaA1Nha1HL+5Si
u2DaFEpxJWMtXQo5QK/rl5q1bH8A6pt73juUA3cpWrfPyGdEunzrBkPjv13+1C+vXoyemHNlS8Qk
xcEBjcjK4DQdi2e8UDN4fj23OOhQ6jEbTCat2rQoMfEGgtkYOzXxjjRWTjzSZ1OXsquclMkNqGNT
2AlFLP6QzxPdSA8TWwooi4Erub8PW1fWVlNJv7uS4JAVLzOYkE3/zAqPpj82u9Iq1R5Bb/9UArAD
7WJjAX+d80LzYU7Gc8GmQb3uZE2bgu2PJcVxeFl0ICUaUsJ/yWXiigG6We3vkB25lA58la5ZNzHF
OLZ10t+jYx8vq/GWQ5YsgF0V3t9ioyypht2b2QblB8AEzoN3piodCXG32BtIoMlSf3vrnJ20Yxyt
z4ByvsJ4hxGVRu+c4B9XblFgCoJuiiicHm9c9MpADeo2C5oazXYcPK4VSgKaLHvmjpTm/5ENX8QM
vxm8nC4awDqZOHEUFrukFsc3NmQgglJ+sX+kaaB/mHS53hjMVMlQW/7fMT5TJH8zQGQGYPnFoPCz
EJ2v1R4D52PFA604bR6sBrB6cCeiYzAk0kc/4St2v5gfigkKpcJvp2ITeNzujsQBhHPRehpve366
StSKAC/2y5hPuvLi8vf6x4kAsGlJK41w99GywR4iynKzmdI6Jeqop+O5UDxQ9lWRcrUpnQxtt1tP
9/+kWfVMnIdohSKu6QDIZhWxW9gZ100OLVr12K3SGFhNmfqewXiFWJkvc/YNXg8vWdBy4+WEnBDu
KJNmhQXoF+rlXFp7wcyMDDlrqyRaCQJVIu1GVL3iy/lwZAuE/idR3lGkSamasZrkFzforwztYuqf
fYvhc0ysc32Gpd8D2NwZlVIn/g2X/N3io/JyuHEEk5ak//9NyMp/dq9W9xuW1+8LnXLezmWEJz3L
ACNbrd6HRLZ55CWb+BA8HgtiZexsNlzDz8bH5P0LItImgzad0tLlAyx//+3FLmVjX/2sUmYc/6f/
+icMAdtqox1DJS+UpGcrrHqOi9cAr2DGT8Q5xYZvXHEGVaX18hVlLu5ZY3qkB/9MrYxyPkXEK2CU
A+sJ1NIxIR7TQqWeQW/OY4k4n4p76KtZ3g9O3wiWJAUOSiIlCcywhsoops1gfVKEVn7myJu45X42
VwNJfztzCb/xoV1vSoEMsSQcCwPQrSxHXfJrBukcgEcCkJhWsLkm+7FYb7oFqM/mGHeUQZkOuKEx
HmoUvCnk0PN70pw5wuRLfGzZkRL7i0KxT93D69Nex2BQlSNjeZ7F7hC5tvYe9Ib5ZXF1DxEOpBA4
ey3RPysy0fRWOv3DC3XqWdWYj0rFDMZJwcWhDQYzAaFFE0/qP1D/lt0zjgSSaLm9DFYhzVmIpr6h
C9s6XlZBPKeWH4hcIM4fQ0kn4DEz2Hzj6BI/LFMeIV26h+btYs8qlPvHgj5FeJcEmk7bzhAZ/bLN
d14X99Xifz8o6CcPXplFc8Uiq0YOMUpwc4tZD/fiUSKKUXEbEQO8qZgs92ErX11KjXq5MuwuPVfL
mKe8jMnzEGLAl8bF5Nx4tnel0XeiJ1LvGURjC3kW00h7BcTnI6e1kYZVCKGFzuBvjpnbnpfcEFRK
kSHA9xnY+EXG2SVLFr+IgLnCymnJulUFYT2eni+Yi6AcxGLXkcapxN3nVsr9xVOKdPNMsmk4JZ7i
2rbTNkaSkgT74EcmGUbkZrBpcaZSMXfc2aQep45DTTZ2hZsCz9vU4gGv73Q/J0tsSpqJ7vOPpXQU
liNOLXz+a4Fdrn+hrHr5kPUW7y2k392RyEwIOgTvqcXngTO1lr7x1lFm8YhBQiLGrAN/oG8Kqa71
2WhZjsW2h6Rbw9/NjeEJ18GeW9W8H0ho+rPn01gX46sDAqbTqsuUwd8CjVtL9zcXpzy7Po1cRajW
aWev0EALgH6gmn1kb+gzHXqvzw+SDbcjnEOEXQq2fj94E2lgWKVc2xbnW2OaPfBVyrQ1UZM1DLnX
PbyJmKz7g42caRiGHnSGx8yIwtOeEuo2EuV+E2A/tLibjeMwBTulXkwl3SIzudAv492RrK5QtCzp
zd3r89jTknW2qBIAU1iptUTuew/L6sJOaWfx2ASzKErQV3B768+l7lKSHubeDdyz2vnp3XEnAEGu
NEqTpfwmW3nWEsimIZhhZdC9Ke17ZGyP55ADzk+jG5HebIqcFrxzSCGrd66YKvvQq114IcbL8zTT
M0OQ2HgsjH+pGe9DOalXhFmPbMEl8Lo00ySQstH5MnzWQtXXbK5kra6Q3Ql7YrfHbmO8gZwgXMwv
EyV51PYhHz5uxuNkQ7AudqgBZT8puRJKzVIZmgkc7qIKbyVARFmfUDHa3moyPysBQYqlDovFcaA6
9xd9Wr8/75S4lfmB2n24dFU6ZkLKBhUrHlwjtnCL66r9WJ1PHnEfSo+b1DyQ9wlqVSrkvHqcFt8B
FfY2yM8A1ZL+7po93noAyK2RTGT1RuALTokxOVOsHpbiQYRTaPrJifKqwcBuNQBs66DDFG7Pci96
KifaDfuW3y6VrJE7trH38P/148XFwXxUsyW/R0rs9Fa9blY4zDEiUbLiFIuxlOvl2B3JkX2PI5lZ
+Rbb4IenhG5paXHsFF0zyns+1S9QT4AVRJqtALKzTuHoKnMlOHiF+SfTBsKBBbRsI3DGUo9YFiYy
MnupYH9m0CavdRVyCHv42q7jTPxTbU5Pvg8ZxXyVTfei6ZZRl2rmsj5A9dxyKjdLUXyYdNx95M/T
uCC15i3dejbRz7NfXi7gsuDRkh35C2KjeU4YMQVVpDm12s84g15iV8/KRzgU3Ske9OWoiG96kSpB
dAvf50tcbqIt3XOR/tUfNuCCFcVhnNRgecBcDVEI8thzD+ZuOosu0tI3BkPCeLdpRlgMsMPa7qiP
FyW7WEzQWwLAeCxOjm1GOlb1JIBtaIahnqVmRNf3o/Ehls5RGqnvXD5k7NByv742I8NAj/ghxXSj
0UF388uGUCjA2tQQ2HVIBlZoGBVw1a9POXhPYtqc1kcM9ZbBfQipMjpmVrgGvC147748dY5gQ3VZ
5Ef3/lQB+YIfyqdn19el1AKEXEeq0LtKSlBWSxDhWVBOQbWRYJz7el0Cx/wZJncXDg+biMQWRyzk
2sUwUb/ZPKhTxDJgLLCXtR/b4fQp2Ogc2zyVmjU9rpbtOJKHMOCYcMJIk1AAHcsk9+A3NLOYbiNy
b1H/q3HlnML3CLptqAn3JawsuYIUo0WyJIAw68cwIDyZi6ecFSKzGecXWhLpwOK5DlE0E0DjXAQy
rWKKpKMAcu4AZPVOYUr5+9W/pVocqMlBcq5HKiw7wkxzSoVsUPURH2AR3i6mahH3PyPVnIYpvF+D
C0varrtjJAq6Y3NLLdWCPTcGcvhY743yS/GMO2cucNh0l0H9hbvTYKN6Q/VuuTvaxSwV4vmVH/Kt
RFOE53rH4itkFD3XckUQDDjmnX/iX7c2XbOAPp46Tn8CqMkqYH95A9r1IeN9hKKnJ8SrSR2SLB3F
mtCSVWA0dIaahu2gbee9TOAxDI+jn3ruGUnmQooDn3Jr+p9UbvIlSKaqhipV3lwyFAMghYSs3qag
XpJ4l0us2p4UueCZvznOJEQeazhSaGkt0jSROzW5DN4xx5a/HWt7a9bSeD4C9R3VIOapYClovs90
MkqormDlS/TWt23m3l5TNHuHIGVnHKNh5oS1hsfC3aQA518AyPzzOW66ZLPnys3QFxa6t6mO3DEx
Y/yxD+ZQsKCDvGxzYcs/Fx+HowvgZch7D3MVVpfezKjMI6H08tcxgQYBHj98X41yRxyJzACgPxEa
ldr+vAYmf8aUy17IN8AJS0h2tB94Y5/Pgc79MwBOLyApg2/BiwQayI/GnM5N0KJa3WW5grgWkn81
XuYiWsegfulMmLAaWdB41GEYfKBKHnk+UJ2pkM0F51/jGAjXp7lKpxqCkptZVq3b+coRNHrtFN1U
mB8kE7Y2MiBfHvXMKJDkMUNB/L2xKdxkhlhbeiOZ2MQhVxxYH7hLY+vZgawEJAJj75w+8zsOhwl1
C8ylz8pI9wIw5uVIorXYmiYurGb3Ge0pdxiSY3CUaENn/QOLCKwj5esNUElY1qbJU5S++JPELTOL
cILb6sIqwB8Vtx5u23d6eabonkJek1FHaMwPq7YCbW6lTZjGuCZhw3sZ3tzShrAbJfCWI2Vr24Ou
wIB5zNPtaVcuT5zhrQMXhUrAh90aF9bM80/oVA9RCceMkjoiAQRKsKFJY9was3u1b0lo/5llDwJ0
My8hFg2zaALwXcbRcdUDylsptXxgzPphCbTJKUou86gV9sJM88MXCZrHPYiyvwMNmv45wGIrXSL/
8iwGhzYxTTKcjwlDGYIyIWdHmguKfCfsH4ZjWwHs/madmJZ2HP6LNRm5+r9OFcj+YCaQu340NHiK
3BjLekZserjZfVDcWUvr7KtyxqtOQ5IezIh00zWN3OP3RR4c2U315hoL3+RP2qkunQTamn9PMA5D
hzMF5esdPM0VKS0l6BDU04yfHJX2+TuLPDSvU8xPLPar5yYCD7oUDEbIMPRsQzfp4DkFwpiAjlee
NANoDaUtzs/axESQpZBVnXh2DUGkRnyZpe5zRojMwBdJsHuxGwXT6Hmeq6RUIN7V02+zJKxnSp52
4JyM3/jrq/0y12ybtWltMgzhSzJ1sonXzpW51Sab7drSKWYmmuAEWdGQLq4Ux255ZJbDLdxevKh3
AqnY/88YNIMph3Q5Sm1PAWoRX8U74rJ5Uyv7ZOyyA/ebGjCNP3F0mMGJR7CTkzxpKJQTM64/FNk7
W/iQapSk4AwQBroYxTxy5B3EQePgEXDjFRMsA/VEQrA31EUPFhdsHd6BiGb5wQ0P8hAAmFW0SE6Z
Hd2IV9qWbIn1TlEKnEht521Ev5E9olvhThl9f3uwGIfbqnP3WoxkFU1lAzvWg2HN3vNBIVKB0Ein
aheCJC2218Ttb8jUdSjJNuVzty+byEkyZ0oDsaMEkPOAYGxq192Tv9KwlA3ccr1Joy0WvW4Qu/MH
hRZjjR69bosBh9WE9Y1Atd0suLuF8i3ZRCxdnDRfQP+aGxIWnQx3P4xrbDNtPp99Nv+5uoFmR6Td
wVnkaCsKxU7CAGW8alTHrwHxAGjAKQXLmWMp2Zsa+gHZxwzh0vkKbbXyGbe5U6BmsZbrE5QoqB9n
e1oVgzSNbX4+hd8HoVlfFWrK2b+u/6RlL/M4Tqu+evg5HCEaUTDumGJR67tf+G45TRxwF2ee2YN3
ajFS8oPEE5Z/M7+Wj2cUMEPSHjVWOb9A5zxrqvaFw3fF7yLTF00H0AsQqlDoAfk6bsY7YU2ma6D4
VwozPwaErs6btTjqinrBXifY+23sgreVaKSCZyGI8/9xPGBonAN0OjRKGvxIVHpKy/Num96MpXlV
s81DJ0iQm/1WQr27qMsWTBT85DW2xEikqo9rbR6DD2UFDgkCXY43akiVcOZXXqTemyXS+9gsZ2zH
bX7rKjH+dDk5+9jgHrWbBcHhuBHC5tE7wqF2Tg74yk5GHzJRJVB/Y1DTHSFeiWj9yqgiuIxLy0gy
dd+2iUnW5F6XYuUAzd+gE6onxGI/m6ZfHBb+Iano90bbMmmzK5qa71Zy8i1ofHjZENQXkl9fkuVT
bR7P39CLSIoEedDh4C54MSQv0f3jr36NjEuwdXvJDURDtL4+Wigy2FNeJmcVxaMsASfuIz0naYTr
MA4UQwpjCLSTmiDMS3pEwPRFhnJaof4MG2S0TmKGfPjMWgEVbD3bGXBZR2GbF6VtLt3Lme3PZpVu
6/bZypk2+zVYHkP3NN4xNswAEVVjWsGz7Gvbcwn113SmPrinn+6HcfSTfAQA/KSArHZBOS9lahJP
xS89lWS/zbl13y3hIpe7TrIjjjzvcMubWK3gKbT1Jh8JtP15zDLo0ifumHkjjO1/psRM84w8Wl7o
rRTQybuH4PoFglPKZZXVKo4N1nBKqgApgAUGDq9fA3l8CPT7zFY3+8TVnyeEnv2ESUoPi8iT1MUf
+jpBq+6zCaNpVOSuZYw0SA/XMwOEZJ4anncwxmEQiTX/zvJ+Rw5poFSLLfZQ01eBXC/va+zL5rj8
w03GB/yhGsaOqaBAvDTd7lvJovS60V2rbqGiT1yhSRFOj3RN54tCRVqKfgNXcMUnW5TrxysnxBMO
Z4NOqyHjzI9njIaqC66Ny2s5izwWT3TbfTjr55nXgvK3UuzYsZpfPmqONHZU5rQ6KdenXroZpOOL
38+3wARGY3B3r4qjE2/qBJRRelwPeq0lOk6kAN08mDnIU3JIA3I7aBKnKJ+8s9CejdEe2J13G8eI
QR98cO4kcnIZrM/XdgE+LZ+ZL95j2BSXqUaw6qRpL6TYnjTYy9pCgmTkzEiaGJkTK+lPH5coY82t
dNknsPMIZRG4LuGNSUXv18QqcaRIHp/F2kW7JyZ/x3yaIXcBcIX+OfvaY2r62XxWkVMDfIAf0Mqu
SI8CDUAmvePTtqgR3CPjbw2gzNhXorX+cBlewDGij0vTicYLQ4vbucpgMaFZzAaph+mCtnTWd40l
8ZSKxbzDjKZAealCUbczrhRGR2FptGu5GynfoG2NOgrRhAYiTuag0FOJ4Gq+t/es5AprCYFE9ju4
VPsBDViO1hqgLULhBThsPlGDuTcWjgh/uAq4129w48fcsqIxfgyMVY0LaURyZZI93RKLg+POpg4/
kP+x36CoinnWoYwPEZXB2jeOgbhjP5uMMAe+5oSHW5chym/fKTRxnAPOGWB4wqdrJ+qsWvnosUDH
kLfrmx/M7NQscn+J7KRW8++ZS0KN+EObaqSOipeWSvr8rv/iwZi+OfUHeEJsAARoR8b68wwjcsbj
aOxV8OThB95EuqhWd6pKHkimZHcdzQ/QBd6aYzsyIFAuCoid4P1W4qzm1D+znY4R/cmNKJevTjt2
JkGA55hoLCnBiEZO7wDXspjO2yZJ8lMl7jWmwt4uBHeOQ5Q0+tEhRfLYyDoeAkQXPDMgRGARlHes
kJvG0FysOmt21aLoiV4LKjOBZD4YOkN4d1nVaJvHwMUIJgWYMhoTlQI12M9ikMbVbFWUpMN/GbB8
XTvJVlfmJN+CQmaU4JL363aENjHqo4TkspX1xG3sKJ1XLyZ9rDwFlh+h7PPTW/w6pUTYuV3vOm17
V0OvC0wzGWh6xtYVfAxmBAcCN3nsdTpyTCMM7z4FJFv6+abqKtiD5Iz/sXjdFuYySQLLkl91InLb
9JBrN5lj+GVo0rEQsSeIaJEkWxZkjhdRxpVrIYdhPiNBFgbFIJNqxtQ7LJgF4btiTDDGAcSB8fIT
3Jsj0aoLSqzJAWy1I6/AZon1hVFZdxj/gE1MpDyx7I1rSL4l+/FUbobw5kfWVaDjqdP9oODLYgNn
gYUbssARpOxyMq83DWvK4DSUYvUQQyPaw5A4V4TlJLBnHu9tPJcj3HTv+wLvaAwFkaZr5NWuhehn
J/m20DsnNKkj17dNVEd3HOivsvXwhjOsfMwLvFexybFitGPliL17jF2bjf4P5LCgGxTNwYU0FK+p
CULuKKjqS/tEKcgPkc3CswUIWK1GkwhQAsYZI51YC4tvs1HxlPPS+S+/yK4dsXculF9potk3DLKJ
VG2uElM/lECDs9LKGMG0UchOf/VgH1BDezoNs8xbsn6BF0TblWSuz4BWukOzxots7gNxmeKVrMB9
0lHwz+vN2wa067ifimQ4vJSFy1zDWH39PK332A8iEyHRpZc1CpAaaFNGmCW5EGu00mQBLpOPzEKE
XbfonO8dYDZmMaBEsLCcxu1hcuQXD7DnPIQjzifjli/5sqMPTkrTvW7jQ++29EtN0yhPxavGXqtA
eqZ6Znt2QFKQef2yvZZj///D8rr0fZ8dud1FYuUg3smuoF7esUbnuTPVyA5vGWnNao4FJKDoZSV7
ld7UdLLWZJLFevGXp+DHp4u/7ZJRvvkykJJeuRz13nmgBiJUpIPxBz6p3VaB3tKfcGolKMJpgzpH
0pRi1Iaiqi/nilUfuZ2yqn+t8prXE82muW/cvX1b5f0dXqITSY8wJQN9XFrpr6e/JhON0103986t
NzhEotyHvWoD8aVJ3aBH7ZhtwULV92s1jeV1TfmvuDbwgA0A9Nr+rJ6wAoAC1z/7vYXqM73BCTkv
hwVa2G/vuKMk7lPBqQMRjB4s6qth5Us9cr6MamxL/fXhdzhVNvxt49EZeq6xA+rMa9EgsBQuPAse
m2D+e7kkFcSPs9BxWvuNqjxRTfdC19mLZSb5hemS0FgWCt9gXPlLkWDRITKxtBcPsD7xhEQaI5Jc
Dpn65Ww5Wecl14J07hUuZ6sD/48A+wl56AOOpJG3K/umrB0As9tM2xpSPEYT90t+OLCrZcve62PV
bDL65luG9F0bhKL3gNzu5pp7Qts5lrYpacDNrQrwdO9//iCzsAz52vXCh/39clcs1BewwEGdEVof
dgibxEmSgiGN9wcwstXN+4vdn+FUuavxxZr+zdGsE23gmrDL/4gw5wojirNF62Np8HosPC1Yb72n
g24YF4UBu4nkpEEze+lZFDodRfpTWFYQOCNiIDnJ9xF2Du7x5INZNxUcB+qnbvsms+wwl2ivXPbv
VjRCliTDUkodSblxYkhs3oGH9U5k9DDwQEO7A/bDyGowzMCWrc6Ugb/2taeIc2A65WGuWck05zDz
t/jGSJKLaH0U4w92cbiqysMRBv5AUwZWB0mC/YKvpFH81HteXflRHzJBvNoyGcNDzqv5A4Rg5ssv
Xgl+v2sQ/QCdqPaJ9eQAR48gUjz2M9Uh8GirtlFNA9curGR2ucbTgkVWt0nzl5K/64CyMz4Bg7T7
/ZNhvripJKi6ygyXPKxyrbBloSiOaVBBhPP7aPPBsanY44eun6JqBSCvv74AfaeHY7T5cWsycJnM
c2ZHKhMXhgtjlF4ZzsEwBt2JMBjPYcHNtBw/VLoEY/C5uHKtVFf0JHcxTEByMCwhYhPROOu6c01p
sB9CBe/aajH2tRT06J1hBIxDlzUjTMJpGKfMJ9tQpRb91F1mi80Ar5YRHi4zjSrE0VO4DBXdTl5a
GG9UxN3a7U65U+DC468gFwdsjQ/GJsdGZ8Th8r+L/x9X/qT5ok6+jn/qwzb09VH/46xYJXaLWYc5
dJAajawx2BHNQvzaJxTZkHTSkybrrgCQkOJhVxb17eSmDTE5QAHdWaIXJVUvVssOzj0lTPWdfgZ+
O/gZQAUgLrjreyXo3XRRA5ZVE8VOUgbw36rsHqpiDkRXt6VM0vy6EzkgAaonXjYFVlYVSlA9IvaT
13kEe4pMtQeVMU0IHm8xPt7JlCqCBlX2hJ0GGp8Mu4uigfa4MPEFkklbFxJyMFDsGEhjLcSNUqUO
4zbNP0PJ83EzLSz5uWlEGJdjAX8KCw+Qj/ze2+MSg6WYrDJPleGGFOXZIEM46oBQ1o3Utavtjk00
PfpUWXNQ+f4JyznIoJrnmafTU2S9NUP5dxQxg4fj6bjtbtvyFshDTnzousRckgCdWDvKnjdneeVG
o/PQW8J/x0NgleAFJ/cO28WrQn2868x7sCU2B0saesS/9hAHL6+ykQp9fGtyzr3PHvbLfl+OOqxL
rVBx/2uvoDGVYCKSwzEaTKFlXrjL1OI8zoT1Rc4iEqLIyiRJbLf/UOAuECYKVj4U+KVsRewSYhVM
m0TiD5DhRJFhZISy5lzJOSbZIpinta93nd03ZWnwr3ASV7Zsp6eAF1krZZw4Vfr+OS95rbVFQoEh
2azqU4VpFlgBClK/b/f7mlAKjlfYC7s1JG/hKJzZ2A77N7MbUDipcqCCNYfo5CSL8k1/o7uz2Aqq
1Om2gNPHbUn3+6qUmbHanTGHGWS1x693Jbr7n0aq1L8zs0/pa3PD4x518J0ZyVM/w8++FqkNRJYn
chev80cYeL6uTGtxUzO1DmsGGm/GRlfqA0V1BmKCVMAohyz8RRMuOk7R4okDcUoMdKljCcq7jLFE
LwAhpbWLDrXVZPYIORz9UOd0Yrz+CAdDs8/Gljgl7ftUkjC8LtGGkeRGMwEa9INO7ZSguPSnMx3r
iHE3ICrroju8hYkU8fydaG8YIV7s7+e0xAA/FfhtDQvZUJSyxCkYjJzxEOuO40EsTVqUzNPcfoEn
ar8XYJB5G4FamQIXCkeSUMY3S/fXZcYFiklaYhvzJFGwLachROzOX5wjZulP5QyUZPpKLJfFaqo6
aSXtJVW8VuAfz2MVOEX4iGmnszhV21z4D2JUv8aNL38PmRKlegztBaBt4EvpNZtwITWQV732sjQW
WhTfc2KpvE6yYScHvCDAYuTRAp4kDHruNiGdIzvAkG7QWUbb4FK5JJKOXYKpa+brQiFCzQ9Gt5EX
AmVIEyZlD/0ePduusdqc5C+NJZAb/U/fUWgBKxGZdZBa39S+SmzXg2pr09M4tUhk1+ThRRZirRbU
BrV0u/EZC/b5ZIfEoFiMtzfqm7LwudDGgQ+SguvnkTpF7HrE0PaWT3LI/0szwsyiQvchU6WqIfQ8
qCe2ZfnSFwsxH2+g7WYBgmLVYWIUkfGyoroZsalljdWAM4ojHtS8Y6Vy/AzEv666tifPp0KDklTY
OBbx/76MXexPd7Z+pDZ7QrNZCCS/b38a7dnLv4tJsgMkBRh1uXWZTpOD72pDPk8sxYEtJ59hqlll
SES2gZZGB1sRa2lznfTObBJu8S66cscIn8GUlR1JEg67HFulCjj+RoOENSxeuKIkOA4fQxM8+/WZ
oaefbXey/UDqZtoNWWKxlbJQDBjQaPNvLA5MotkqK+xavoOvCRiQKGnDQdoo8QC84qhFQIb1R2C8
FWK1zUoFH1WMjr/AiARe1P6tMnBC9KmJba2DwFQnUK5rhlnhEdfgu0DtPbhubVYoj9ekcq49Zrq0
Ara1lsfy2aOpH1KvlSbYHWiwJsKxpk3zem5XunKMZ2DReBkfmI3RspjWGpLqUC6ucr5iVOVUXSfc
Uw2t1as0JwvpXvsFU42y+dAKQLOe3gkf1CLZz2LOBbNRqG1iRr7QewbvP8ICGeSpQnXTKfWDgfUp
hlzeAhrfZn2WdR1P5yJd5zOAIdftyL5bBIcXTkFKr6tlZlpmeOScTec65k0ScPB/nNzrkY9RQDZq
msW3W7JY0dIYNWS01uoO9dFy9hrbRb952uPpTTrrY/lSbW8WSXFQjcBxs/B31ahLhZxJP8r9QrYm
7fij1dDJ9RZLtKtJm8OmoZ/RLCbNGm+pZ7XjpWObs1JuvRKUT5WbMgAouqAiqCmP29Wuad4P+1GU
Z3wnUHztN4VubpdjzfrV32iUMKQ43J6CvxykMSQ+qAfyBBXM0uvcVpYzViHuaSYFTzFU7fPjE1Y+
S83TjUFWXyplziPfibmJJ35/OzRMYwHfQ7v77Jq4Yw0OtOGXJkus7tGx+o4VbbRJaoSYPWn/fzHe
dZQ28UAU/152P4u5JBLZ/yJLosOj4XAWqSxhc5jVXAqmrRaC+oSjfuD6sXDeVqtCQRtcA8b90ezg
Qry46yS9nJSQyRyO8gytPeTXF4sIKIKXWQx6BevU5l/xvTgRVfo/7gbJosBHSW+NsgFhqPOE0fo3
RdQbjlzdngGehS+NjYsspyXdNsxY5IBMyz/8OGtE2+zDN8cug15lFmkD2HYL7VAH64R2AVxngBt3
HqCPmykemo4m0D+ARDUsK17jG5S6Q9tPO/nekN5I9y/WjyKTLoXzHciZ3/cHVNPAE3vjgpfMZPTI
2XINWaxhvAcFmTZl4op/FPhonUFRAUIVHKf/oVr7R2Z7yRayvCdrFBhfwqcJQadLqqK50tBLwVrm
5+8Eut7j60BKyTKtpK3M7V/VtOtnaGg3hO4pSYkfPqtRin8Zm5Cd7tker5Io2Pk3IAWSHDF5JxQ3
lrODdA55kry8M4XFq0InPWC026gyw5Ffg60uxi4l6fx1rbvUJB4L+YMvpPcpaTM6Ty7DenANwYCq
ofJ30qh+KHhwGfPWpDLdMztdk69lOD2lDfnH9ezsP4Hu6MD6qhWE/lWOI95h0KoZWKb6gIgUIMnR
d7bybXn7PoCfxq7X+vtMQ6gYPgAtoxluyc7RKeGAMhDUL0brMoTMz5j3VkZDnfjv4iXczvffxfJn
ME0UV0pM4q7pqkG8COfBi6TEBIuhXi08uHwZuZEeCNEbyIU8T3AwuDHfpCf8nwCgpiXhqxTFV+2e
P330jRrkrNGS6cNXIjsO0vA7p/TF40/Cn6WgLo1WrMyVht+OGeNxjEGLFYxhz+eRM75OHY59a5Yt
QHFvZPFVaS18HYHj9CJIq2inR7lwyTpkgOl1r5Jl/ddLFVOLUFXnwLKPhulmznctWsyVti4k7UUD
gOf86YHu20nljdtjp4XfNT7FDVsLrENsioWuH+LAZNaySAuvU84getcBhqJLsq3haHD1ZgyZnJXh
dJH/gwlh5sh+nESQm/CTFHbTUrhWTuZQ5SIghQieH5+GO1mdvc3x+DrZTmicTYFxvLI6KBo6C7li
K3cFQzjgHyetLe9smWOPy7eZABkHCf3V1IKCx2LJiFBf9VQh/run59kwaWSYE6rW7YnIXOobQAxO
teeLmce6W7pyAUcv5yJkLJSho0Ss8KfqnKoGhSUq5af1fmhHsPCLlTomR3871LbDGm4UOoJ/8CIj
XW+bLK926ozWs+euDtZXGikIYuB+ykZ5pxVBYSiuz7TG8IbH43G4bUL8Par4bEn9trhHDi3iXDTv
MO3bY0YEpjPjsOklzUY11vSz7CqgzFeWLIZRtD7GUnEOHW6qXjTwEmOaVFrRMTG9t5UlKhNP1EfL
Z7EMwfhjoe94kkTSWuSoXgWXuuDYh21kwvb4lW0kJkq9Kx/+wWl2e/ZL529ez+Bi/U9TSNkElE9F
YJJTrscIPaQuJFdKCTSs3Jci0HTlTtS2OUPePsJE96XTkJ6ta+riP8BCzs7rVuk5yuRTXDaE944A
Lh1KUxNkuo1nWZIEXHDmTpHszx0sdCUJ+xXZpo+XSU74K+oscghDSjGbZ/F4qLyJPcTwmdbW8NLm
HFfZU79u/hVRGeZXjbfCy1hiFTP56sgvagTDrJ7h1mzUMKBCqiYxdFAQ990o5hLSETPW8yyioAKq
IGC+yv8b+fxHkSqFSjMnjRcl91cqQamoi+9GHaSFfQY+MkkZj0ihvXPL5GxOh7Nzb6TIHd4IHcQV
n3K2lg1QV3+eWbbzmLEiVT4TwTZt24lLMmLppYfWegRzrkbtHjonsDInEwHkHQjSprq4DfvmKC0X
oC5VY3N02GBywBAcJLnngS+KklB9DIQ3kav7ZKKcqagk0xsafCt56fVNaCCyXF9qjBQlBye154lW
G/+Vm/5fJcctFngzmBUX+cnhYFXycwzHo+FkYR6RZazIYzRGlHsf/Sh1p9IHRUtw7PEsAf/M8xPL
IgJknQk1RSUHudqsc6h8lc9bJZlUkEPhOfxWM9fxrvOTNblTOJT/Fp5dTKCYrkGB68fDDzBZk4tB
nWYqlAWFrGoDRM95BiZcSgvIpuXW8WouPnAK0lXdofiQyN/whOHRO0AmbJiWBd0oHuxSAdKjXsm7
jXDPFgL9hsxS3exbNqlgZiPkhRIQTlK+0vKntHCTy4zNFAWILQPyig+zSdDcJuF9hQcUbPk/VY49
oTH2tS5AFDl7HbPMWc7M0U2AKwaOsbhp38Ped7Gy8/ODpric0qegAYwL8L9MoA7Bohzkvx/D06PZ
4TQImjinlBcZ+ZIvX/w+At5QubNQzQnyck/KWE/XMvfz2mb1CNUyhp9kiBIAoIurXcIBPHdMrBKg
8cYYE/+JzyZ6aH4dtc4TSr8ZhfPzFNeM9FkFxK1x3QVpjYq/TKpzBrxWKIJbky+PIFmVb7K7ZAN7
jUa54Rk6tUf2cdm87N5e+a22RYFg+7xENlykmx1aMuHfnNX/vH5uqNP2tyffLqW/KCtt4lx7vLqu
eaFA+bpeA5cf6yPDsn67jWuN0LybdIeL3B+g/IYbGxtV9/iUoQD1OhQ2nWEhRa2doVFl1WFifG0c
DKVLaV3DZXVkkQF90EBJYkZmTa2NNkCctwxuksBOibf1SrPQE1p4eAT+M+HrUbskv0LexVa1Qj9O
cbPx0+yCvd/nTW1DFH7QTuwe2VozYGo0Y2YB8NFs6lXiJK766iMQax++GlJDB3ZK0IXQBZzIwD6g
GnCrh9pFmAFlSDq0Lb6/1mbcmrdqv/2LHOHaF9mtJH3NYUofAf6LPJ9VWKK5o6bxu7aE7bFcC0LI
u7+k1K/SbdouhyJGuzZ4FX5W6MOxBpCwBSg4dhde+5cUoAkdCb4AtVfUMmbBK1dTiSn15dDecYRm
8u5wVchYNgSqC1RbQnLMp+EgQs1lO5YSYWlmSZZ6p0QLPSa2NB91CtEEn+BIBtMJ/qa9o4GASsIt
YR8GRFOd6yCPFwz9KU8+xD7roKZn1cRyCJfpNhcRWsiPqC66vjY0FrmgMfMWInTy3GdH8uV9YbCf
1Y5ZZPqb4vOmZ66KcGcPrgxMrxerfs6VGxmyzK8ROb+owzOdELSon/UE/VWZKEU0r8eZ5nXQFGIO
lKYj8tgOOTiK+sxTqpVm+1jW0eyAksDXJFvGW4pmzzfKblDkAqeMktTG3b5jHSzAi0lQBrQbWEaj
uK10ZfODP6ffRO6DYdJHAGWc4m4PK0wyZa1XVNHvumDSQbIaVx0rPmF+5eMCfIXGZRTxTGPu0ceQ
Vu1A3CuNwdXCc5dm1U5vHHFCP3Iww7GBb7ih1xeQZCqe7zKy2G8g+u1SZpnZrZaKRcIIlPUyoLk3
0vMIJYw8Ss/AydXPqFVPzRVGriU8WDGItyggjG8e9NokgosPrcP/Dr6FJ+qxKseeADHkzOBu+Xie
6nrJL2st67I2Y6g2j3VR9Gp/LPfBByasiPZdSyukCoANxI96g3bPhL1hDQ5yNpgRuugQ2GWKL2d8
2D+P+kTkkkgWKCM0GQ9a94NwpGX+8vupUEX54YbOLEg995+OG1qRrndc4xyvFb/OPjaw3bTXXtXO
fCU3e334UGgjBCZ2pD+CjreclBQQwIaLPf4yPT6qB6gBMyiPBU5HNySIrX6fMcumY+Z7L/aDHY7P
Us9hT9KA60J5Rbq9x9Y92BU5aemvzCdHpDsTtLNrar8m+uBfLYnSrJx1KzZ0bIi/8jWo2oP3vJNf
b6AJr6DYgaqrYtL1DLNEZNbwviEr9I3FVLNOFsEyH+WI59VtDos5ByUwTAjXbe993NOYBifDnqrg
9RI3sonmVfKK/Wd6nHjXMDgFUnYCa35KtupbZTn0csPztOwXdHIOg30G1eqBIKbtt6uhp6taYPW2
ZlVaPK+FDTWatgqIt9DWMWYRIeLAlvJ4OBiQMzDvI6Qz3/CV4Cdu/5XofBI3Z2LDRBlLfq+GUEl0
eSUSc4CuUCvRtpwB7jzknMwRnBdK8kJ5xPIvMhv9QS7GXlkwCpKr/tdBu9/Hyf2Y0ylxFmcf7rp8
QDebsdFjamd+4BhPzt1dvBF3YlW2QxRSNxkKHL5KyhSoyMO/zFFCdfwcBSCfxKwSQQw40cSi4IrF
qY9Fp31ikUwWnqnfMXgVMj/QbuvV5p6y4MGynIkvz0HhLDcCeqneOaTrm1KXNoU/Ji4u29X8w/Sj
MsruRsPcEJFUPrzBUCDK5ZBn6KaQ3RprfmE6hA8M77WoPD8w8qVwCcXgHqYGHliHqfmZXbmHrfN/
jsZ9evLSikz4qLowc2PX6V9yK3WPQWPC3+My+4x3RdRZRWykIXtsl+wLLInjjWDoETZEE9K5CXnX
e5c5jm5dBUyZqg2KzSnHw/Au5Bd1kBmweX+IJmgS6uXRw6xCt+KGJbHBNwjphYCdLScciSi1qR+D
Vmi41FM/zuxpmRsxRRpGZbDyopN3nJ/PdI0lf/e5ENaas3xCAV2rCNpUK47kQHsU+FkLqaykZ24t
3Q5VrYzGgpWJttdl4rP8GkQpklj15H1Y+J7qSS+0j7b5GEGmQrUiME8gQg1lNrC0HdYjUEOYlB6l
f6KrDwzxBpDh7l4fXFLLgpHxDQ5CjzXotHyBKImNv9T4KMPBU3sz15KVsmtAwAWDnyiF+lCuSpHq
WmoOldr1ZQ6NnzQN4k/1vhnme7Dysr5eKea+T6dmw+HJ1ljXjsxsyy2fRsKqLt/Ns4F7kF5dyE2Q
m5BxJlJ0XKFgFI0WwnNvSIc8z0oPxj+qMN31SPIE9MHT6LRkB/lZTSE9bnsuRlqzXLi58gmjC/2a
64NVfty6uel0f+QnRly+aD49fBBoulpc1eNJQoqq94V15W49WIHnV6v5L46+0FBHAALUg0MdEyYG
pe1ewhuk4TxXrr1ZL6wscHnxEMRnLHwLtnHELcs6kmTEN0OZYtorm3v3EgQCTl45WkFk9rUFsdHe
JpKTibKhWf+Jqy6rG8xGD1q+qgYpM7rwibSP5e+12ldN/birRkrK+euGqjMiakT+ZOwFZeDGDSZu
gctWOGqrsfFGthIMv3/hg3U2WmL8KLpulo2oGpG6hbmEaVTAHF2HbMThn1tPjJwcq9pkQt8BuBWP
490/ZKwZtVTsknSaFt8iCNk2WtMj3N8wOxRCmVGzmvjvCvvvojYbpqIuQU8Irx/i52s+HnB5nnNO
74HDEXq+Uf99lTQbZ/0glMRTgSXa+CKugJtf5cPlSH31+g3ivAuheThwPs8+4m85D+pl+wyqVIlW
UV0g/hCG7lmHtnfaNTXoTN6Q0Ypw7AXnb8JDNmsnZBYKTTppIBLQIdd9iJHDcGotiF95ndaVLpxx
Si6wD0h4/Crny3Exm/LUZGZhYUDFJHcL1EqyoMxhyTP8qJOYyfmLfwYMUe9/TCU9VwpEeNPl/Z5T
AJPEriB8t/B7G6h1cwBCJ18p8IRuygDFIXq8WRDpcIQqyRtAr6paTxWVuhgzrSLI+/Il/UppNpyU
ap+oa3dcrVVhqxjuvZFZbXfgrZifTXbUoQlneEplYzJ7fuNIVtwAIx1alqYk2n1DYgxKw5T4EzKJ
hfe+X5YErd05+cdsH5daNbI1L6wF+P87dvfzwPB59zWXuZizU+NLyctuG2w206EK8baXHJUsH1qy
1NEE4Ii5T1Te1NzoX7No3kKM8of73fAKzD77rEgp2GJB/b7WMIaq58qh98sObAFurmMESTwmZxOs
GG8vl7UlDbar7e9O8lWtD+ZVLxInTOMz/UD7aVb0DNkLZMjNainD1E1leEJ8qucTpmzvY7cZibaC
cQQULo4UUQKF/ktXv/zDPElG4WgWOf4WBjyr3/VmlxIyykcFRRHtK0NWUO03F8aOdJPeP1EFLeY9
TY702yfWzXn5/9Ku4/ZNshVRy/1n58Lqe/lr4FdMZPdfwRZ8WooV/nC4bCJQsPmx22MLsWAgh0Xd
7CoylNqx+qbLslAGaSMGZLVn5qz+gc8QdrrnbVlAc66l4CeoR21/4gMiMaiOobXF+JV3X4J60zSp
l8ZLv/G8Zx1uEZdH29CPVPeSUCtlvPvUViHoigAb2IFgg79/NINXDOP3BXmHGEp9DTMBJyKBEQzw
vpoYuIEheQWKzPPmGoytPfpf9gXIApv9g9B+1VAb26nm1U9FcJZKmkeqcXz1m224+/8JItNMnCZ9
Yy3J4OmcN0m3xM27Pm4zVXTpoJTkSexO0Bzb91cUZuLokj9S6YabAiu/lpKK1suRAXDqBzYsQlH4
yScWbhdZdOYbB3q4eEixMPRbrXLGwzci6q+XLGA9lEGUo2XHBKw3t8wc4Ovq+oCWTk3jKmlsHn5s
TL3sZwzO++Wc6s9zd/oJugUqHqUL1toTWkyJhIw6aGMhwHr9FdGldY0JjCv2Z4TSP31pyBsFCnIn
T/Gt0TykpFfFwcjfcTHLolo9+0seJwkynohYOOPLOjgOkQ7GQLKZsqswomQFccSXiALqHRjPdyLs
8Nfre+ILgeQS+p68SeLhsrcDdGs8unWht3zPW/zYcVfg4P1I7haIf8c0xbcnHsQJ4CTUMntAPeJL
xs+69Cm+9qH4AUxCbm3vcrphhqsbL0hMBe5UtwCmhF7n9KvaQMABeEB5VCN0bxfPKj+K1s3OWpsY
xIf7Nu3wOwE8genIDHfaxUxM8TH0bTf3ME+QAl9gyk1OHYmv/acZs/MM6/W4oL7GC3hI6xv+8gMb
RtWyApHiB27iok8wPDvLVIqoWuphvf56p298KJx1tN6UWvN/qP8HJLeJqfi8RH+HxkPB8j/uawD9
cfS1QvSX/6N4EDjRiK7kVl5IwG0U2BF/2f42o4GZG6jK147v9Qvqsl6hYBMIb1eGNxoY+pOPZOeQ
KsPEuHorTaLuEZQs+CH3AF3Mny+mvVuZNM+F702KvTdvfaWBCk8hLQIHD7csqZ+MOwtb6ZhpMF1U
K5AMfsALJ41WMZoknJEkcaiVtR9UIKqJZkvl6kNe4ssG6nyypg53UKMVWScXWmEUj7LV6hxvaRuM
6xS4MbgNzEDWF6KUxCDI/B+8mzks7UXkaKf9nFoj4SuCjYenAIyfCkI1Qvos52+GQKUxsjw79ov+
D6Ox63fJDSpl21tK6269RtmX1rBet5s2vMW3288f73HBgud4xNKQhAWU/4z+2F6oQj5drehNGn8g
64pBuu1dnFz2OAKEmoE08jBY8saOujyhYVvhjnKAYYyKFQKKmRm1HCktX2qw+xa4JW6cDGL5La0G
qzKi9CuJTQgkRk2Surxnvg4SZrFHu/3/116SqSuSVCJStZa9r15xdJTsi1aWGlQLd5XJYrJUjuey
YN8wcuN+vmhQUsGFafXnSx1vYWO4WMjLnlI72uj5ZGCF3cKdiCCqpY5Q+9ifkqQ00Knt5Uy8X2VV
WnGd27MbJGIUPDx+QwHh1PWBlSJ7YS1bnP31+ATpZOD7jZnFg2qsyspJZrBJFlp0lM4TeUy0vRov
sYEHEepwkotlfXGt//ezig4F2wA5Wru0CRon2Hw+vp7iqztszMf6hhDEZYChPh7rnp/kDJ5GGxzp
36810N8jlCSOVK8BKjwG7Fjd0ylyAPbpcYhRyycGggJZEG2PCyKT0zs7E3j6Ha3uI37ecdr///Ax
umLR3tHVTvGRPEHvcM9q/KhJ1PPc9Vc6Vsh0APxf3IWNoLO7HHn/EbWS88J5oc+O1R2Vy16PlSbE
+Q377bLgpmoTmeVXjLxpsxyjtoulDsPSIbf9emolgh4JCvj4z9OoycuGspdMrcC3yT+SYqN3ocUA
Nxfc5cd3NbX+MDOTPIhZwrBn8KSgTIhcSr4UUn+/Q+P/6rv1na4yfTVkKPTvB3IlY8xE50DsyF7F
igCnbIBo++9rb0T/nIoKRcZrGfW9496/paf0Hl6GjykPjRpNiD8H1L8BTcF6BWZ1K05lj+BcZxUT
9UX70ShqUFgTi2kB8kj0Q8o2M4FCMM7qIrUUmpZ/i7UnO0/CjdonxmTiD3rnZRMcbfK6tIvY2lNj
6ppqbq3X20IURYKeiiU7nYSHhb47nr6lLhGBOAIpCdCe8lCwCNmyhgJU7DVZ4z4XZEHXoAbHmQ6c
KVlMmVrvCMLGD5QVT09UMYDJ8z9/5gdeuJF6uaSZCaQhe10oFcn4cPe1m0h0i0EFf3GoFNTxzsGE
3ylfHMzlUp/g+4tCZQfFJU1SDs130kPlq9s9SQz6FfLr/zQjhqxNqcnq/XGyw21VVVqiM464BTyU
riTQdkMgyVUoCOmNDLVj26fp3mXPGFI5hOi075ipxyxHkK5azUdpzCRWspjOxhryK1avqKdBESx1
4PbusufTjr9nHFhsVlGk5PHUlvM7CTENwFuQEgctGQ+Uom/nXzHVtRpuviFPBY+s/XCREzbPPG/t
JuZUj6ghO3Y4beL9L5LqyYbtZ7rQdgSMdgz2PHW2URkPz0A+XWz5y7qjhTI80VHgc2soy/XK0syL
JcOHDQKD0J2AWIIleoMfFcrrRfiAeAlEUQJ7BaC9aHcWUZhD9/SiuN7N7wmxN4bwtXIKhQIKZIet
h2jkbyY8zftQ6jyn1Swy4pKjVz0SavLRfK0PqLpuSqBAKhP6zRUlN+bOQ5cRCSQgBvfVuc2m28to
Sn5urTHDgWgHBHWDKNK/1N+FXIQhyiXhkytrWZCKqkEHneqsrWBq3qEKgH+bWZWzWKkNBWbor2Ip
S8AykzipFDz5djXoqPmiMdKMwYooVxCWYVZE2Hmrc2q7K3QHZhJrc7MhNrwVG8QzJEL2Dimyo+He
B9OckRxodADZ2sCfRGNzU/rqnJG5zZ31BHcDSOrA0e7MYO/Y2oGE5lPwP/PL5fQXcjBQf6M+MGDy
qrTeo09lOaAOYeZ0wMaqLg7sBf8zpOvZdr9z1hk4RPuDlZNmCHfxv02jY3ytitX2gAkOYE/+oeX4
PKb29105mFIb0D06+gVvOzJZEfEs5BqV45jKiJqjfWpe+gXJF7UFpmw2oQERQmfJP+F4XU6TIyQP
RRS4E6NTSijXkU+JzylfTYvvDSzLVfmokDRE5H5S6D1VilngclONPsNcEwuLA9EzIaJxJRozsLko
luwWaHK2FxEwEFGPT2AaHakuon+Oe+X2K/MWd4GldX6obzBM9BjYbXYwDowTh+lik/mFKmQ+NZFs
4Zv+G26gF+SHgGGkOY38ZY8REQb8+iPn7Z4WVxMK5iNSYWAwvOnHoNVbWqyhA7kOnpG/h1JLnliG
KB4VfVMVFpqd9HO/6YRyeRTBNloJKtYKEdtKi+VGoibrYfsUOF24CL0FdNH4671AFfr31Tu+iQe/
WdLR0Qs6U0mG7fBmbrc5HY1leg2WKzAxJgzF/6U/US4XXc1S+Y+hQW82IWCIUvkFPuJGfHjeSyNN
LHkrPFRcbm1D03yY3L2sGAaQrElBj4soa1T1bwiuW0VNZnJ//prezhL8GqEaP4W68/5ABBSJWKEO
bQWyd/9IMlm2EDxG6GLTIlPtfVgtQRk9NcgCGsIln4ui/wWHCofh/IFKFGlxqNH3nT9B/mV7mq+X
oHIMKJZlh/SB4Spzg72svFmtfw/zOlidtFEvoctSPwqcPOHDx+CTgeWbkiETy5YxOkyeyIDTaYba
fJCmhrvqSYOYtgFPPG0+lLXBPmEn2OY2T8EuE6q7MHYeSNceNucOgMcp+zYE32vqWUQvdOY1fr1m
gboNTQ/sL+TujOrR6jN06B3BoWpX+hHQEOGteVtj6IAYZAfN+lvWzI0Iw0gWUIUBxiMRbvMi5o6L
g3PB/g9WV5eFyH4wZ0cIcnJ6RX/sXxArIeC5EWTIn0BTTUxxEzVtu0ZD0VpnorrMQxPKoVSKAOEg
ZtIbo9JXkf0nJaRR4szW45BoB7iZWgMn7B4lumhariF1uRTnlWHLG464vZb0ct2Z70nd3omiKMW0
Y8FXk/ef1Td4mruBLvWp8KlBaerewy9GyktBR1nsEZGzSdLpNO1I9SLhhfCZ3i18jOYJedpqu6Vj
Z39Z9PObN6LyRykhxLzxpIC2oj39sC7Po3cQG9TDJLa6bnnePlZG2BBlIjnTb3vMk3giUAjs8Xza
R9zmPGpCN743ogNNqRza+7Q2AlpiGrCVC3qqZpp2mcI+2uZDPq/0YGXSsGg0XJ9QHvNofgqPI01u
gT8ziMr8vo9DyGWWNlpC2WMnf0mkbRb/nkIQLK6K/hT/WzAXL2yaUnMcHyZ/s1p/AZS1Lc5DXgP5
HBsju9QBKfSP0ZXFmtPf3XoTHoI+zStoD2KJKeeaP00YbcPOWnLXKD6Xj3cp7ZKmi2WXn3A45d3S
JH82AkCuPzf9PJgrSzFYnbyYNHSOXwRfAZp4IOwb3MGCD4ftT5qbDcoXxBPbYQQLmGa83ifSUGYx
mFdd23i182tRe207NWd/KZ4KaiNghwK8/UnADN5ErOalCV80P85OTCHcaIZhi71eHfIoXWv4AP59
Il8f0bupGHzckKWwNalOEVV/TCT62Z7ZwYmcmc54gmFwYxZovY0ZuuvRFXEa3bAwE2es1YYpN3V0
YSsIZz1OYGS0TkzpsJQuHa7xvapcrJlZvw3+VdBU+SFLrCObPcqn0gENDW7SKbvve5zbcNs8BZOJ
3xdezjsjZTcJlJQwsN1SnsOnDQtz0B0NZZS/IamY5YND+Dvk4E7pGqmnoRUYitl4lthu284Jalie
MvoAQbJNskMnpdcDck+Nr1GtFKHH2rUIl5svCyNUBCq05LQy97/uUND+TRAqWzFZcxicODZlq5xn
LWb+hg6F/t7jEdaE7VKmI2yjGjTVnivLeGsM6LvfIBu1JkTEEJMkIKCbhHMACi4aUFn8/68ala72
6EBv3CQb1rCN/vWvG1I29SCjiAqDWyPryaLvTiRdOVcsx6Z3HvwBH67oKXoFmsxdBpdvKuSAW4Nd
3ZRZM1ItITnHcu0Rzq5ZVb3t9mQ/J5NSvMwfOyeoCny8Sx1A1DJcY5E+/GZYU/L4OEe6pP3wPZZg
BYrt8jHGuwc57wJ0tH2PMqdr9aXHj8XHJplmY8XBe3j39k+T1HHW0Dz7YEq+FoNc64fU0yRklSrU
yNx3fqF93wFb3N7EnuW7CY3icQ+ZUJq3Vraum5+bU8CUw54JhsxslI75inKKUnJlIMwXRwqnYrME
HRo1D3QfsjZUsCFrk31k5ZujTRHaXnyWlEXF7O3QZbkw2OlUUdme8yvWVtlMDzEWZv+sp/TZ0ktH
nYyRudYt5f1fHAl/8LGt7rC79snMaA3VUdfFIKHDifmKKqR0OyeEEPtYzHEwJ78q9GzZgdWoa6Ea
u8muvx+cBEWalp9tUskWl7qA9vEZ5lIfTCmQEB0pbAIqj6gxJrJXZ8W1JvxMhlVNthUFit2Bdbgb
h7BVaOFBRgwLJrgilK0Chg9UsWVqm3IgkHC9ghDl5EHx9cCVkVxpxzSM9hGe1zBMxo4sBqvv7ezG
Z20LStnTDcTaClsxSHbw95hz3A/ybaRppy8WV9XFXV1e2PDbCkA7ygFyWNcjakSBJAijIEBDutUW
FJbrFsRtmXMwAQOyvsNcOkhFq7OBC3dpxWK/9y04LZ/qnMkvZAO2Kk5Y243YrAFQsNKD6ISzUpmx
vxfrxZ+UBCXeqBuZC5eKiP31PySy5oETyTM/pVBY3VtaYIequU9rJYa5Ej/sCHRCGzWRiT8wjNfe
GAIv6xlBWYibIdbqiW0vaBLzr0PQSmxRkqyeu0mtVujnOcaDgEIMr5i8oYYQZXI8L44VTHpxzRbI
xccluJDREEH1mDcyC89YOzgzFX/Y3cVvm6nNrSikEBAOajR8p+XVyhtaGbtmBAL4DOcfZyRlM7o1
NPKnOiXkbpVJH9XgpuheQ6N7zYHrudXPvnQc7CiLc53thBv+yizSBwPK8ONQ2Eq70niGc/J4jBPJ
KCZVs0tmRPc6qj/eLDawk6+byCujhk/CE4ue4gcjOnR89sOxVjjvniD8J2XXcGCH1MkP4W5Xon7n
GREdwnzZ68YVIb8w0rzSPoj66on7wA9dXJ1Nu19FocJd4kwiYy7CPzMnNXZUiQfCSJd9Y9fiB4lK
p8L6glUnab+zn6QZLClANtF6UcIfARnsFN/plVIYAdH4z9mXDJ3LVJbHe6AtadnsIPzFVd1mjv2p
ilya5/1VfDhsQNlVAL7W7evKGKBzTSctjlOWzi8yaflkr7POmdb14bC2lczHxqPTkqXB7o4Y+8w4
vDS5j9nKEC7Re7rnvMW8PgHPg8yZFg22+k2VwQwXssM+VfdLEzj58l/E25iJ236oje9z6c6HQ7A+
f6FWwKCX61j8GFFq/5vl8fnywHwtI0w9aV7SLtu94BH10yyGjyUh0VBCGbRTLv/iGapsUEMDve4Y
5jLq7sILEqJgcqRVgxO1kluJvtmGqbCCQdKZ6o6oqPJqB/rd2RQxWHinSMLql1vL3Fr0nGjulHAq
TA1D5qBAjdRw7k2QnejOua0uQWhDvounaFKfEcAcJH5c9WXRyLMg9uE2cXH+ox+IgsBE2TTgvUyF
Srkuf8cs/HhmZvwzjkCcqgsQFLfLEBKAXsxl4guSspSiZGaGxoauyNMWAKWzBLIZbIRG678ZUv1g
fEcOaiGRkM6INxuFUr3q2hYkFW//oifKtQuvXnRKFqHIceZjsqsnJhrv8bM4StN8F8HJlXrPamfb
kgQelMJnVbNm85km9KhmOwL9QRVbo+gQ5KFDQ2wC9k6fw3GnFYx7tyZibmCqxEgSFE7gg353VuVR
ZjyrvZvRk0zp1RXl26l3jhjvXeYeLLy07VNE7vsMJHCQJvbXKZNsGVl/nxsWf2McWh4Yw0QQWHKf
7RArzUWd3ul8eF6EYCdumpYO7EnKMaN222rkHs4iDJSDrgWm8wfZ7NikWhkVRC9y3ssypbfYhxBT
MC9FAzUoakyUZE/p0VaJuk9diQmrkr/oOm8IWqa3sNKKPswCfFFE7IT+V3fhD7oihm/yU2srK6cH
gTC+Xnew1XssZMfA5mH/17YozjJAB/Ben/pufN5J7lJVhgvnOzDkfqyLJY8tCLH/frvCyGqmeiMj
b84YMGdolwbZqdkhoqsR6jg1SPIpaKD0r9LVSCalvJFDtzSpxOHaZqkdFjlVMj245FCMDwvu4r7e
L5CbOv/GeEAz7O46w0gZSIh08AQN1sXB10S6o1SLP1qSB8vl9jELSjLdqhtlOD1yi2TifWqYsauR
fkSMk8iXQnAgfZV28KWxpacaPAHa70CoOzR3ago+odR0cERQnVtdHRNfSw+JFWuC+oRuAFfXrV8C
6imZW/6/gJHuQJfBMGD5wuAW273UoEOVjDexyUMlxRjkzLfdizYXXHkypSG/Yc8CbyAZ3dT4t7W/
SH/Yle2jw9oto7s+DUkVoAvci1tthDIcMx7OJt4bB7iCMq3BeS0rC2MMrcFZSwHm70WVY/dObOS+
DTkTI8Cg9VUEFsv0RBRW31psaMSIoqOGoL9A7v1dMw0TwcU2gM17UN4qDKuSr8iM4R7/eVUOtk1p
7LOXn+XqMnvi2BAkSaY6yl8aAcy5KSnEf+K4E1xKMe8D/M+VqlJE+Z2Prufm4AsNt6lG6xxTJ3Zk
Czbez0QqJX3YV1ohssdbGy0YUdwDoKajr9pQXT4kX1NwxI7xcbUI0Cju+rw0NHIa/K1ROWRjizS3
qVG4vhtFMH4zNznwyCAYeLyhDTPBgLs5L+uT1n7JDBMESDOQYnzIMNwLptWum8xvXmP6FxDq07E/
r5KzCZoJs0hYYNCiSuETK16DVGXxco6xASpXhRcjbkjW3QMQ51UsPuBhtXVvUVxxQ9uCAwkLoMIZ
QZgU3Tyl40TMPpPZ4GPh5qoEk4RKM5o5Fb3Dyl4TYDo1xMlJiGiRxAvNJ3CfvBtkvOxlhnv/7gb8
Val1l9c4+TF2Gp1ZVAZS1jxhWdDq41hSy7UDTFMm0+ba7xIzRHv6+qlwxKjbLqO7Gl8WMYQEUmBg
IBaMqZUtWaMNachBvR9sJ38WLRyWw0mfDJkBdeYa5qVQPcPJpRstQolcbxG9JNfkdHblriU53HJD
4GR3HtWyITS87wuWdFWN3SvJcWn6KNE5ZRk0zi1fkeEnypfx5g2fvae4omZt5KL5k3ghAcGrM3gR
PuTei9x15TAAN8hSYCCab+k4kNoi0G+53dkl4KPoZeVZSdkC5dowGxIVQzok7L6/JzFJerOUHC3n
cy8ZDeIP5kqDIemDiobvY6QL3CUuZwHFXTEHvOupE3YvLryEy31GccKgX3b0poIxGpRP/xPtLB/o
WmviJB4UyJkvxmwoxYUH+TXfXzBEaLcpbXcbxmMFKpoRtihUF9nU9YXiPt22EyUpwASwjuJSaQgt
ck2tVpA3F+Tuw27O9nuW/jHrUWgF/YruTqY51998CLOY1TTTwL5fCZCahCHPUzRYBGOiIB70SWem
7mDnfReRSO42Cw6NtJY8/7wUrP4db+644aioE5ZCaUJ0zIl3NvOsRYY2XlXbu1LHkypAhYrEXaSz
ACirddNG32zLMCUovEIWs+27ph1DwgCYxq+VUqNXtewyFmRS54wcVywfuPg1ma+B/o9PzCeKyD3l
KHlijUMMvdLopLnPRetH/fNZsJrkY0KM/9Ypcn6bMykUO/8KhkBhNn4aPYyZCgbio2cEtiuR15k3
lKLzjYiXYwUxp8qk50ta+D/FxtilPYyAhptY3ArcWYaxKBST9hYrHEzA8MkgV0La3y2WSNrfqkOQ
7QGc/ABNm5H/XWKWvCsrKvld00iFf+v3lWqek3OdWkHqzlWYDNJg0NK5lwdwC9c18aNvsy/aEJ4P
4nK7v4Pf0YJ1IBdmJGzHdvlkeXD+TCxkx9akponCE1eB+a8rfo7ghPkrFSD+SCSft+Eat1pTG3kX
3CSIvoJu3Y88lDGkz8RJCdRfsMWWDtmiZc9H4dkporMu5J8z+r21Bt7HxmIS6oWTZV2UbyvOVs+K
tAKBIXTDlS57odUaM4vy1jKq/8CHjFfqzxFw6mHO3VlBB5/8FJH/qGZY8XKloRDk0DeQLETJntAa
98Kkj62V6xKAJvmYG1yl5jKamsl4NbjxXGHfSt1ci5S0QiQ/0FH4sloQxZZW/xWrY5wJsD5EvfhO
0w92tYrTLP6NG7ppE+qZ23EN2dty+WwC7O3NWsY5KhuxYrSmpqJVN7/DoA09eKYD+AK8o6sIL3y2
df+8KJDqhvA++9hbxVVY73xiOkrYZn8m/+J2bmzHvp+3yrX14C4uQxJMA1wHGbkvQxOdnBCt+vxs
HtsLhvim53Afr3EA7yOR9AfgU5eenX0namG1vPbdbBxpMNzqVGTK0f9GZ/fIAN6Iiaea+YFi86aE
LwzaOtsOuPwhtJ4PVAyoA+mOjruklGqOmHcexpualj58xC/UGKbonm7JQKtwfe6pVev3oZfAIGGR
5+KgckK/ggU/2ucuGpUy/x6ZrySewWstg0Vx2MLzAipzDFllRgcHPm2GuPjt2HZPRzLLrA42q0vA
PW0bhATC+8A+U/PLEksqi8pWykGYhlrglhSWeClXOFfUGkODc7Nw7nR0tFLtrk8BW/6dKQftjBbL
eIBvfqxbm3rRoDXvaDi6iX1KckwnADHheUUXLwAde7YqHdEdCZT9hBE4nBNOs6KAIedb3ceMAKia
L+SlTeoOV5CvviubKXTeKyNlyJr1sDkvLRS2mU8FCTzhTbMUKv4fVxInJ6Iuznp3BNUt9paqhB2o
JCJLGePh9/Do/FaeOTNHbE74u0iw6gvyfMIfkqzN0p9gHigwtYuJdTf5h0Cy6zzESqNN/gnODuRG
rW2GG5NJo/pgGuEvr8uK9DfloQe8fnYvt7GEo6VpgkdIAdl7kuLVeaBmYzCzdX4Ye04tRVY6sGcB
OUPzqOSTxmKPyVq6kgr3595YJr6nLRcZI/K91X3VA3diZEvb1A+oOG5r3fZxpfoOl2dMsTnTuIBw
fBfNqQu9rXaL35MAAJUY9lbPGUYGMr8hruO6xzS3wW5r4c5+GD80LLHPhIk6sr24nNeX4ggEMwNY
/moHc4CzWugPVpaQu2AnyN/hUPe0feKRBMMsGbZ+bEXWYaRYFXTlq0Bfd2vq6869VWrOh9zTSbUH
hFvJ8YClGxPwe5QRENH/UEuIjRs/JgeKrn2T0tx53W3sDf9ke25WZ8J8KyYrASnShuS8iN4HbB7S
ueuwRFERuh28ILk2nMxZaiWP9PPLhn8lofCRyLlYNvd52fbm0YwkUov7wEWi5HbPyqQDwSw8jnZ9
N0uHwV9trcMRs7vheSVgpwbhSvsrzVPuEaRVHfMdGw5Uq+zcOaWyfN7e8zFPwX0cVyc+IheC9RWH
BnMnDIiD/dSrLoo/otp/0DkEMt3iJPs3mmttYfi/09o08Wops/eByB0vLMAMjnLeEAvUK9oPISNh
ls3kQ5TKZpgFMal7+iSer/EELcF6/ks/866XuE19baFeEvfWQOCY8cqqHlUBjfO1AGiOD9jzRJoh
ck85UzCw57YVLJj9kJqSu1/BU9DB2D45Y2V3ch9cbzN0/kUitBA9/7VGcBaFlpoXJ5aAZYgRpE10
H9q1LxgHFMlimF1ep3WI7IU1faAHvzChElIsr4jnCisrg/yCuitZH5wTeIubtDv6H0CdxLF2nVLf
Jy7iQMXzLYpEvADgC8odZLv4afr9TdYfQ7wAU2ACRGHM87baRpo7U5pYUGchFwkv4J9vFTW8RiMY
/ESOaqU5+/PcHKsiYW83x7dUWuDbEWomqbTXJl2b8NHr7lyK7DPK4xfkz64nt2GzXcjSOLHZ3FgO
bUe5xqwbkA1Gy9ja1Zpn2/QFdZGkrA//I6KcPnt2JR4ml4/Osk2f8+baPU1wP5uuUy16YwiVQVzv
c3cfIKCh4xssWoBb87gtnMXWqm9FRuZelLGlpTBFtuLqQg+S2XMIIOxw+MrcfZxLc36LNA58Iqi1
2W/NbeUmEf8S0lFXokOLNEyNCyU1FSmu58npIJQVWZKgHIGW9Tgyw9KgOjRtu1ahiJ6Ca/1tlpgc
7+SC5d+iaBr73p/YcDs8lMG9FH0622LlFebaS0WX1fCLy+54MacFDpTlj9ifj0E1s8cSayELjtTA
j6/xASh3ykoSULb41LddwEHheNv6hQikv8LEOLouUfMTsaROOpOqBNIgJ215jYsNugiXg0o2pWsp
XJAttATN5yyi/tZxiA/DM+KVIOOzEs9flZBuaWYggU0kD+toqW1RsquNn7brESTDWU8fiXrRuTLO
yj2FtfEkqiV99ePLwwmd22JIQCiR6KFrofaf5MnxFKBp1yHCcIDpjf/+lYuVuhGstS7RAmgfwV4O
SZwL3YgqgxnPTXiUMohuOAuZUglxyO+DgWpVx3C9IhsfwVWXZI6K1MURP5MvVBXaIMzt/ZFu086n
c/4TOmvG42hsHlV9/2L1Kl6LZDi4WwDkXu3gDCDwCr8/c3LdW/7xnAwIws+0yRrmYc9F7mrLcIW+
J3CPbADt6xjwaqFFELOVMtxHB1oddk0z5YhLrFvEWPLte61c8f+MFOfv0eaTUxxrWMLPYlWBUYXm
O6GwQVlDhn5ArNHw8C8U7zoy2EOnQx0ZnEU3Cht4acoYLeKlyBhu9S75BxYIbTBsSdrPegzU106v
ACYSWuUJ9JBkw6rW6ysxWUu2N9EsMGz3ReTr/uDICgLvhmqitdpcgJRJbuJFK/gp/RX98TxTQ5+k
dXaipDX5wkX5ZrLRm0ML3IKgsXQ2z5V8G1cT9miFYY0PqSc7Ax+pkWHv6uAPFT3B3/g6NHeZrsmb
LmXQeRDiJVDRvngBMOF462h7TjnXoLMY41L+tAZz/tl3Dp5SKUHV8tGUlUOTTES7S/A2zGAFT49O
uaGkimtp/dbNlRdushuuvmHy85kAyp6S78S2ROgV9SgBtGglx3lELOrEcXy3b8AiZPPPinCdFc4M
gyg+I17kDRC02mePHvsJqBYK9p0Nk5fJBCG/aKfJ9F+u2yOENKIhcA8yDuNwz068Bh8T3JEPjdta
X/7LK5sAt0uh14rN5u6Vjpldl4ekUwa75Fc2Wz+uwuxjqRZJkr3qq09UiTOvUtSTk9lXUCZ9oovL
3/8jrw9STcJKw+pfsGDaQS386UBUpwCDAfzMA4i4d9qoLcJObszYkbiWJYKKjQxZQkr65vrM6rVs
KXfyMyUVlQK++ihnen3/VlXt3lUPd7PurOldcaY5GPrOgiKcflaoAJ+hF8qd9AWzCt5VghSD43Ic
SztXhz/EoNFa3d4OPeycyiMrcGt1Diabdy32iZb1ddWGkJCG0+GeOTP1tPJDPGy1zrKLHcMf3Hfl
ZbKdAgWpgyiEN00hb3y0kRBbybCXQETrzEmfV8XLvIufAMXvkG65FsLd+PRenN9cRqG5WywP9bWn
+cs2Kl7Bt/NlukNgVXCMjweng24WFBm3PiZ5JpF+BSshir7g+jyqm+wiN5MKkpCVE+YfSl/J8Ss4
53jsYMOwqZ045lrfTpOfwQukvKL4UCOeRegbhsC6pVsr4AWZFRL2UYCEOz1UHyqy1dMQ1GzagF1G
19MKs2RW9dKzIavFFvQM5OHMuc8I4pmGDbYYMcv1vjXoiWtI0SHzKSeIq2J2SQ854BPHN7RH5vS1
4a4uijtaEvAEMQXj1A8/PUoVJmQiYe3A6xx0PNcrb4Y9uwtuTNVTyKvSVy39LSoffhpi7HunyBjI
dIqy0Aygi0wvmw2A4lRmzJz7fWGRSpS36a9Z4Q81q6D8RtFduj561vQae/2yrGaOpO5dfmvtNjxp
6G7UhAnJ0iOwRUZ75rOMp766DSgowMAU4sbr2DgPbf34KXACZ/prlvhmHfU5ABbnJsx9WeyX+Nli
JbH4EkmG2FR8/G/EjGcztF/OleNWTlEsfWTUXFtRz91cNXrxsjkFd3VwoAS68PkCpH8FplaSWzZs
2KR1t5fmFcmrKHoGAgsIFxj6ZJNnDAiCDUwPM/2AxT1+hExPhHbmk01WWpZIWkPQSYw6Vmm6Ed05
ORzx3nF1tTDcok1yUu6dyCfWRfqX7daJc2UONLZfQ7pdtIcIXqpy4d6SAgu0xYm3NlspJqYybnPT
lO8DuBzsbC4hD8Y97d8l6kuIDzpbit2fKPHgwZpWwGIG6gidRHXgYtFrbUQYzINAQnj6SjPMIwXL
CVPjc5zC5H4/GDzYY0iBb+RgxnGHy1Mynu7PLyiLFLNjwhz7DYNRKGHl2F9f7CtVY/Zk4S9vduvd
dTg+T49DTT2U4r1mLKZ1Dl3ftIVexvMEuv18M4qxl2fWGoUxFbuwxgs+CkVkWI47de97lk300UKe
bFHZJ44a9GHLOquVBlpKynrGNh6F1dZ+Bcq3mZjDPZVCJ9nE4MUj+yvSuZTuZn4F2tvP6I2bhEjJ
O+uYT20wK12baZd++088PhS7/SNp2CdfSlqZh+wk6Cfcqn15GcP33Y4EqUj5TycrGMZyEI7VNDaY
H+A3LeQM+G7adRWE3nSqRSQqrejyjz4WEADAbAMp/nG7qZlHl+9zZQzYCqeC0GxLEffeBFEg+Ihs
iSxUuRBcGGdjNKTIYZOQ7qscdIPYtze2q0PZu97okmAdpSen09ObiqQGVzbpswHv54r4P1A1IMA2
aQv2q/Xj3htF753uSawacZ0WA0pJsjMgYvvI+tEKB5dQWyvDDts9O2CdJpil1jM2xpsxZraUeWJw
be7WHRR8Y4Ia2bcnZwmsNEXXdge9SOXNw62Ch5BKqztGC03Jj5wwqfGsBJpm0wDeObElDxRM53H1
nMsxzPbmguzhMeVaqd7EAELqJe72F2Y0mldU2sf7z6Cf2tIZU9HHQ1B29XHlGoAcncRXEXug9CiN
1zyZOc39TCOev0iMxYtDUGuLNKYTpSuzF+mpQbzGxZFG/199CDeg01kHWUfELwXedDWDcRjr76iB
3JXLufRmxCvp5UjCeaTEP+D4qJ/FRQvyM7s6hzHSpMpuFVcUh6Vxl74T1jFBYcG2GOyy/cpuWpvm
CZIQxY2KlZ4hXDZPLQVhL+YF/IaBnpEwk/oHvnVzBf+SLi86XxOTt6NweStzeQZIiKdf2cpWfIhx
YOfgLMYfsteuvehuZmRAkD2esvgbkUMJYGkgCuJCj6QN3mekOikN7M764kBCuV72MZ6Etc7V36Y6
V7SIwKImJmHI+2GtueHZPDJqtve9/bKhOfmrNb0mubj1uBtEz3s7BqrYBqYqSbbAYXX64vc1/m35
oAgaJNbXXHOWgA00riBxGgtpMPMqQpElFck3708IVL9MQkpJO/AIhZD48+GohTr+qlnG6vZDjqcy
bj0SW2CugK7AUt9O2Z/D4puPaaGRV3oLYHXKZE8c2P2uL1s1lHUzmX+63DVu83fBlRiof/M4aXN5
g9mzW9VPctPVWC0yOifXNevU7wOio8ccFwhQitzm6MyVNWc6Ua2fCKXl1QAR/m1/H7M6nmFhOOIn
oU+EkR2lOvWVtPZ60PmI3epgnlqgCaCwpN5pG5h2XA4ahhJvX4HC0P119pCRWeCtW65XI80SNYgq
CJDCy8h1hLPQDlr0/nNepnp8qqMxjrfcLAwryP598sm/N6u4ItIW6A2t0SpWeTyCFhyr2PFDqDlh
SxbLXlDI4bROQO+9C2TcdFMXEPFrL5VDNI5k78kc5MhDAsF7TFNhbynpR/2fJL+oqbhoo6AgruPR
QBQPYGejFHxeKz3JcggU2inb1MZEEOHvN0Svk2XdmnDfn2ZogQAOxKe9nTyNTtXpbviE1k/3Opf3
JM9ornNfcYj4vsNiJD3hOoyMAKsuQ74yXqzDwcssrC0FJVQG1gBErnpPxOqW3oQ3kuDC2NWi6zFN
QvyCYzYbR0/VEUVjArYSPqaELdsqkzgjGLMGuqP45fXRteP7WNc2k1HVoM5k5bgeOayZ2BD5saUM
FeqtAFlXYTTuVrFxioqiKKatpp1tLW7WWqBdIWL8158fAGq52SlFqL5n9vghG5qMp4AgQf3+RRmz
0I9AYjhIaQDmKWoWYhg6i4Vv9dXABR6fx6PxAd7M0X5oyXJffua5Sd/G+4bmDN9g/h0HNqEH6or0
9y8wNFOYsscRIIX81d3OrtOW96CCJOUQd4QvedRZgicG/q6oHimeq81GSV0ct6hcBF/laQpiyZe5
t7EeABbZqYDgS8YGWydYhM/a8FsQ8WDW2lJhf5o+N9oc7BrhCtMfdnMo3ydLUY9Zo5WWdRc6XDiw
xPp0UyRP/JaVyKZuh4B6f/+sd/jqOxVqNiuLHiK9zR6JzxZldYIQwcJuCKl8puq5B5C5QfOGEK30
umRyWqN59K83P2bnDbM82f3UbQ8hlizHLLQ8nuZSkz9VFCgX9H/EYRpwdii+DPif4goVCmVJ5Nmz
cJnp+GaLDm9BrK2S2gG7Jv01qF5RmmkK8hLDSLN+Aj2ys6CCplIlT2677AgtO3cMvF9XF+sgvYfZ
lPz+BFibwETXHs1CLuQVBinPFOQPM3nWPL9jGOFEcvSp0jVU9gidOr9spSHdu26Z8CajHZThc68h
8QoU6cM8YIkPB/l3TMZqIPaJvdklqnEuqdw4EGtHDhlc/ChRkCU9WuZI+aOkWN5aPnqD4cxuEbbC
U6zWsnZ3ar3WPCsaTy22IQ8KSHRdNWrii8fQSp7s41YhDePrg+vTnoTxp9kwQB8sA5s0nFYPHbYj
DSHif40RoTGKKhDDt5yGl2bA+0QAYMMe5P+H/LWoenXHdfmYnvdqTYIPRLevNpDuNgomEecC+wGq
uJLGLm/oFG5z63KcouWdGPq2uIa3+jp1vJsPyGYZt+2PiQK8+PQNSSt5+Q+XsDUe5JEFOuxc9U/A
g2/wdBY2gUZ4otfVAd0J/+q3XsgLbJfQHW2RzWpZfYgUQDehPub+iDebtlu/haTpECcFLTJ7ikSK
apKa7jVh/K3VzVhspYpJXWSQ9zdHl9oj6BpFoY90Rj4hcNJxyABqmMz6a8ilFheSAPVrum0UTKCF
5Kqq68ODbPcEr5HFK85e2HpK+fIvU8gIj3PAhNAoleeWZ08nOUZl06a06aiYKIF1+IFWXnMu/0Xl
4LJ0aVXeGTnNzeuDyK1vZAxuWOZbMWx8hCqA5Nueyes4wXpLt6ldebeYB5IuueQdhsnFqVwBFhlC
BTg7MGqgq9WObxKBJhGuHHLbmVpm7jxmuAfwtPTxBbh6lCNk7h0e+5TmcEL6Huhro70oofX6fGtu
KStlVerG4TbR/gf8YwR4372TYVLyZ0ovbvjivLzCAo+yaOM95knKrLffUXAXD8D6IfPdINh6Jixq
L+pK0FUOYsHPLWftev2nl7+qhgQYdjbdzwqy301CzN6T7VGFTCXfUYPfDLko+09X5MfVdKenXYLi
1ruzlbE5vWXyaKctvieMvp0bbUFbUR5rkp0DpdsYMPgYa0ksKpX711OpRH2k9Nt5HgxirCA04Yvf
CUhRP7xjhE1D/gmSED+tJ/7Ec5CDa45lrhjv54gNvwbtXdQeaIleadTGGOTVINrNu9pGSkGFBbMY
MMZ/zvGo1msnUl4gVZaNJ+we+mFlPAM3RoYA8e9rNet2/sCo4/B/I65uoBROkV12YS9ap8hH9Gu8
w1islpXCmDyKpPtPd8hw5jXOohm/E+NhJGlx6HmDbgECBBjtDy6L1pw4NlNl/PBFMtZLVkf1CG8d
Fkj/cPNg9zCklK5qRouotQKTjgiEMnSsGqCqhSc9FvxPSAjsRcVl7mM9BRf1HRiTODz4ngXm3SZQ
yxkXSIobQsBjU3bQlSBMi1l5V2liRGPG9TDJ9ooL0MSYOufL8AdEHB2zR3i9DYOyh0P+owCDFA0e
8+TbQJGZsyaPF0vWvwuZnpAM9JEPLtoNPQPkDaCmlNKsFaTjZBFgGL0250OBRz/2iQP9z2XFIRD1
ZGmk3AGWyUiSEOB9dr8Miw9uSBWQMTZGj54Wn/n0v0HukVoNltSes+XTx0jRboEnQY+VR8TnbQDK
mLRu3DwmHxrxuILgwKs2E/MKGmDv+ATzYOeEIrTPafuFvEY0qMBtLJGL+kwukNUnQ7xbFYS8bAVH
BN0SA6DYZY7sGSa5GKbCYnXBYqk/ren3p8yq7gksqGAF3HQVvdUKszP9T9zbR3/u2Whg0JYZeXnn
CbL99ddSH0Q8zRLfDfwOIKigwc6hz+Gne23Tu57VrMm9iu52vAdvwhmd90eHlyr8lM/Rjlk62qFY
jRt5J1XUBCCMsaUJh3o5UtIXz80rNG+QNiaWydLGTb+Ik3hZPgIoRAkjrD6WFVZcFALzKIbWDfQ9
7L4wiGAcQtLtfkXm+PWBQe6wEXEAHwwLypAQtNtiQ6gHeX6xP0ZUJ6MS5w27LKG0OZLoS19cvYtG
dj0KsCupFK4zi23g6VCpAnkI6hJkvsg1jbBJ+UjBO0GKhaNpDecv5E/M1PZ6nZTmDSLcqw3GgX+v
PhC0KYoiY2PVoZCBVrCINWOJOZhNzNYOJuxsJPqahHRpoylLQwW0NOiHHSpn4X19w+QJ2bTve2Is
eSLU2amzCBxme4w4VUkI83Sow2PEvORFblqvenn0UqjZu5ugOYqNjZXBf1RSmjnbc05pkadeP4ow
cWDrP+9j6LYHUPqf46Xun0UtMJNqDtxVLdtiVx45NDLYRbyI3mKGhAa3AcFhQh3PM89CGrY+tBKv
JnfdxO3YYGBfpIsNuSaZrX4eXwNJklFMo1f1vvJul9IoE8jUkt1/F6RSVWvlvRnA8Qa3qyMVBZ1I
vWSrRw+s3xwycvpd6/c2+oQa3HaFYbFgsILlSvLCQGowU+WJugCOBniZWWweXZ9aXelzaldVNbAG
e+OZsYZCsEZxnRztXXOskw7w+/G05gXnadE8v9QrngkYIndaFQO/1VPcAvfBDJm/nJG9khQIhjLw
NkR32LjRJpwRo/pKyn63AUCh64ItU90JBGNSH0z3nhcvb/kZ2zy9p0ULDeQ2U1gHFrRDfo5FSLZ9
GKjwYQN9UnmHTYI0Xw51K+megoyyaFhZ9yEYxugtnEczrMod7MwqP+1MOWC/5KRPL3m4F/IiP1q4
L9cxHixciHJrcXkG9MzUg/uyOlkOSjjgxdaPvdNOWkdG4ZLSnCvB6hnc24jfgl/SiRJL9+gtit8E
KhulI3Y/3w/qtCH1+gDxYjSRsOUWj/E+T5g0wLAgSJqT/wsXPPVSpxqqZibpNcj6S9zkDr/zfQ8/
TzV9NZMYMGOD+K954ie1jfo87WVHLmXqfSL9rRfvdbk5jwJAnDwtZRCKht/SPgM8XoKXI0CXzkn7
RYoNfUDW5SscKj31RRZ4c4dNIVcew9oyyJfyTRv65sqVp/A/UMR6yzj2bx+SE9uVanYjybg1lHYp
cPaspIBF0caaUFS0fN0IAdadQtJUo04wTwLGcNQ46A5BkBqUfHg5yA6ZSCoBaKtqzQE5P2bbP+Yy
f87oGFxUvU33hnALJ0zd9j8VEv3/dOwPKh5Rq+BLivMsgfcYFa2wShu3Dcto2+yq9JrYblc14VfG
F3UR7wlLC/iCq167Gh5eaY0bHpTzNjYiPh9I2/x9HqoWW/I4LI4bBe2hOpxEZT+aeCMLygHL7XvU
Zwkf5PM7B3PS+RzJNQE6glItT7g9U2KJJnMEwbynGdO/KWGbhDNHoTh8Kqyuu5SgbOhybf8aDiF2
ZWUQ2feriIyms02wdNdgrbKYtTSP9OsFm1ZmtAROZhL9Zbp9gc53RxJNCloDDWsBBhyJWI3POX9P
j0cb9X0+BpllerT73eOF4oncPx7Xr8QlQxOj9VjsBGWRJZud8hxsonjLiBG6TYTa6BNE7VTKV27N
j/w0mPKNd1aIsiKY5YmkLPQrC53qKb5KnpBOFuG5t4+qctuYXxda6T6wVvwPE53VgjCWl4c50ZLR
3r/JDFpY7V9Ko9KfFevdWImQeLyh4o8aBwJIEWCkmvlIc0t9hutEHcjU95yWZRMH4Vo3LUJh0sz4
gIuIfgMS6IWuoj2/WbPp3lMH6fx6lXNT6M7utzDI2QyAmuKL/qrAHZWvpb2uATWzZmEd1Bu0bbSb
GzTB3d5J2D9mbtPF0iP9Cu8oKeW9XLLeu5b7Lsuaao3/C2Pm7RBkgc6n27dLG1CIYKzsMXKHwblD
LtoXGWL2e1wuGbOpLJ5URBNaDTZ8/+pISJ2ZxZbYWzTy23013ZbjXsMsaW2xg/shylLdOfnUq8SW
XJQeoj0siktGTypBUL8QrNQlxycegFt9e4zRoYC3iqxoMj+pfwJgBvStpYdhXXtzZN70jC1au/uS
IX8+JbCjf1rfvEVJxtnCRnEA66Goe4B6gBYAR8IohRbgxkJyAdXV2cwd7K3DEP6PndMTL3RA7FvT
pSN741SyRmd9RZB5WiWpYwwgLSrKC5BGWu86iGA3xPj2/L1bRzz8ZNcQDjXFDbHy1NrXd8cChrsb
cyFT8AtHIy43EclwdFu9qUq4UoWm2nrxgC+qVeUGP8sRTC3DqxXyyqdgVMCxqVd3M6Gpw966X+6a
8gmxNEFuoG2RXtqL6u4DhBGEBUcSsy/ws0+iQVtx/HKTcPBryXg/t2Y8xmvr1LQoTLSTgQ8AH7a6
0TB1fc33jz6VEAYZ0qcxahxpEA8qKLpyBbT6Q2szgtIhv37ojD36ZLvI7VVb4Ukxs8KRVxUkfviv
oFUD+MhjYJxvASSWzn2rHh971vWOuTne+NjDSuj0MGMSxxL7VF57sW35JfneoJjxjZb9K7BSppzJ
YWBzsawC+9BjV80QRQpzuMqZwKqzTTyWdmCYEwv3Qyywl8zV5/WzI07QfsM+BnH+mQRxeW8g/WtF
jL8O+yqbi//lxJjYc033v3cXHnLJDIa6Zmp14NysJYSwibVKqcwOSlALBaeD75wewh9uvnkmoeUB
RkqD5TnyGw4j/ULCv0hh8Do8ok7jaFugRe6lVIFjayUGGTk5zRMiLrtdsxH29wvTz8LB5W+FpV/v
yWVBaiLrnEjltdgIQeK3RsPs9rZGN5/Sz4DeOGBATgP6CiVwXCkPY8BnveQTMGkAxOxEsrguxmkv
Ky9qhhTmB9bwLR9gi1JeKvBlH0txU6V0nWRPq9yINzM24f7x7sQqJODmbgIkZ9DPyiM0XdzmTXGL
f+EhBgc4YGwggrkHos8AjEJ9KAYB2GmSYQILcjKNeaNMGvHscJ0F+vqYrRjfK2jINlouNi0rsLce
HlziACIYJYe1aj0Baek6xLyy8H3uhdtHpYBnJJdrf8bHfe0EPh/b9ZPgA0r7PSj6b73EuiYBihvh
Yx7xggVYdrq7wI6WZ3dp6pRcpfd5Nt18xvhRNUFN/qROEWSDe+j/VJeG3SPZF5QMFxgMjOk2YKyQ
7rhL+bW7NJNoWHvWl2Fa2qedG31zt44PgzEP9vLTB3WmsGq6Z7U9aoAWq9U26TaRa4lI85WY8UFr
mD/Byf2oXp78l21oj9t6G3Aay6l93oFvNlmgrBg+XRINYLv/DoGRUyM27+/qwaiGFWSO2LGfK1AC
Q4VeXC+lltSsUGBAWT+edcTLhjVIJLYLmm58ZUcjQ80J1yRIYxOUCPVGZnWMrIOzBiBYJ8Bwn/Sb
u0pa8d4iGA59JCSxJdLWcyDC4gVXa9bhl7vgf8Qfb8I3u/RapjMNNYQ/fefSB2Eu7/mrykY7iGXS
nrm+2iny/zt8AxGwaL4iPQYo+IikT74shl5uz8ZIqkxVQAanbd8SMf3G6bT3RSEH1yp87+mMKQ0/
VGHawiJ6tyzv2FhydQFlCS76xmmKyt/zsG3u1NjJYk1/Y4AcR11rp0immeSmAs9Uaa/aPdzzKvQl
oOgt+C7fBbQezWaYo+tWRfUJvLrUCwem4iBTfGH+LBV34flQwjeauxkXb9wvq3Tds7TdYCD5BIxF
/MGvvaN2C5j2tqXX4PgXQyhP2IYLAPijSJFF3cN+GM7kpYYyd3M5Lt3/A2tPr//QP9zQMsGmvDr6
FqkLGvRag8GQ4lZbOT3pvKegPFsUophqbuuK1T8NfUu/b11HhzAyZnnwZN0IiY976VFZx8OQVRgn
MS0LvrwAvvthtY0zYmkP57VkptkhBQFn3wkpIiJSb0lONCX0Ho2w/0OGn+X7/2DX7KMxYC2CA3+z
fRwJjwdPNLOaYgfyY7RRncQDlfKgdZFqXlkwBv9RbCYjr9yjQFSMMC+b5+SrxRJwH+NoZYUEhYXz
M76moJW2QAIS7V8JFEvXSfEy49toOPpylE40iriMEu/plOTh7Dn3ZwPsasbzzrO5qpI3yzH4WTlN
H2OMBALmOVa9CWZeWMFjshkR6boTkHch5sxpAClLnANYbhHU6XybXsoyPb7qBiL/E/gJ36+OBbMU
gH389F73OTfxQxgZG37PNo7GrKaTfwGreWShe21i5GU6glaE6QuyguxrU7DJYQbBb9T2gaIaAKDT
xjUSGhc49bsVqWwrQk3pWYu2rw8G9ZPewlfWPxFtOx2paRJO0/SRR7U7ApZ/uMpffZAXolwLWqrs
T2r05CzjvSo2W7UBp0xWMimcfWckaZx0hQJqsT94i+2ze0v5sswxSC/n/Lul8PxAz9FXxPvzUdHm
zXFEKsV0daQAT/R5TKEdib5F9ItMa3ezMRYl3rWKZL97LngKL/4o6/ZkEnIK8Sn4nsv7922VWqyN
VAXB1cRqorrQ4J7318g3QtQIJXo6n/ReHgsGc4AO0HgzFRPDvJgt5X0URyJM1NJ9Hmj0s2gWwHb5
/OmoOAPp3uOuKpxoJKS3bZhaD2aw3AICdgd6+uXPqFVFgII89uBqx918diFkLdlboa5JDIla1rc1
ogyA9fJdPoz3VsFYDv1Fdyj4ut0ZnsN9dD/3KjQRtXN6bvY91p2iK8Qz1ziJUWjyxziVEfyceEKm
rSmuO12SE6dEnfIGVjqqJWu/of7NVii41euuLpLpF5bnAGkTAbdHpM3HFgK6w4cvdSsPV4uZwj4e
yOcur6y2W1Nz1Mrfc1fGBj74aVfNqlq+T+aZBvyImrrCdBdu6z6jPXiwJjoi0gTtg6VX3vh6WYx+
Ejk7oRKGXuZhgt88ulYN2P2+ZAvcAw6nua+ti9zDsX3gd8FT4C93Z+a95ZmMIvExAlApS63q18jP
WrURVNpTTSm85gIqc3CJH/J0ZpbfsCGx80G9nOmYkY0SsjtBc3Vqx+JRRppNlfCmIWnJ2Itcp8si
c/KTaug/cQe5+94OEEgagKSkvWktfxp07OZbmoQe7TEPQeFHi4vUlNv9R3d7wlup+XhoCBPbhIn8
fc8nSkydOO3tBGE9UhrCkVNdL5zGQBcbWkLDKoq8xeKTkQKWtAjP2xfpSUZtkI/k/K9o78Kkt9Kf
99DjB6zYbUv542zRGLDYl/zytjOLAUD38o4IWNsxnXPIx+0Kg77qY2/RgmY4cGxVkuX57KvoOGQa
dP8JsV43S4+cDOf45NunhnJipN4tSoxec36Ztt2fgqUlGWvxWVHbtnpkyntFMYsXMUUlcbosvJfe
AsSL3boCx70UnKh+iOGahxRcb4vCZG3jrNKcasCtf6QWWSqxoN7npK5AC52gcUsrAyFch5C802o9
ySGifIu1NsNWX/t/s8o1EKLpWCXMM/o1ICNlPFo4fQJos9DQxa68UanEU2oeUhWOwWk9pPGy6KOS
41gBBtwrStqhkmXc3o7dcK9e7Imru4vQOgREJ8gCgs9emUOaEsKc7cYm7CaK1mLVe0SBkFVBaiik
0Qr3XRKICLXs1OfgiampZ8a7s8le2JElA2piHx8P7S+Z3U6kZ4oaJ3aPbFNOTatCeWFVkzzDsid6
IPc62U9fdHad5xuw7A6/cv0TrTltAiAVAntI9SWMnWHOY9cFujONOjeLa5dC+j2AazTmpidKuFa5
qLw0i5oV9/qtRPyxFisRVyYIMVnZ/kQ44UN0jChuDRIQo/Mu9zvTvywDq5QvKFr0CLnDGhn6v84n
3dNDJpZdcDHXE4YGjS6+aPzvwxHgtFNxONP5CfLH2ejQSJuF5RdppXMJzAR/IsPtdXjEyZCf4T0y
/WRwJwfeSzlrSUl/KQSzkGr85G7HIbiwbSi+/b/P8MvTV3RU8gctbj3LRpzjCVVQI4iDXq4Z/qdw
mjtiB0r5J7SwUb/C+xTU/ZV/qvHWxRlyeZDrPAJcnfbXam97kD7/1UpGCXTqVi6GWVZfsztYhQNI
l9jXqRraaGwWgI9IpcdfK7oeoii7wSgj0zq+IBgar7M3AJO5MigHIZOpXno6lTUGyyk8CcauLBO3
szIVoMyuBKWncGdWN0dIHhqqaZM4CjUjf8VaLJ/8fTvzBjt3P5Wl3iXR8AjiZ3hSIEdgvLmn+M7V
Tvro8itL3rccjGyi9R9OyZT4JeUpbgg5SQIVEL2q48RAVJvgtXRA/oocnS+XQ0wTqPpms/9a+uzb
/kvuaAJgodMN5ShfGN+bIT/DOxVTIGSI8QPVt1GUk8zOmVWEcnm6J+JzpN+4Sfwu3TaGlIs2dNNi
9W88hLYGXQG/eS0QVETpRkdoMnz2Buy9HG3qbuYPor+PnSF411a5g4wu9KoSm8tfyHW+jzdwcm4m
Lt5Z2UmixBDCimUGuGziLm60AtmehIUAW8RwlILkNmq+Kd09JAPw5n4s7oz7MS2k8IsjvjC2sYIX
HCpGVkTXiOVNXxEpOYXLH3wlPbqlXKWMO5DqqB5y+eDK2elSyZlmlHkvNhAm8fxOapNdfosOy/7o
40JF+5WTaQL8/b/C0cgiTF+qPOP9f4dOFLdoo5PKldjtB5bixW3o/J/T/sc44vOaH1PmdNfLLkv6
wQcdwDTZNM0CUqB5xRPrNWhI8VmvwLUYAYwN6aCugSlRQSKlbU43ncyOo6I8GfVB9lBK6RhApzfZ
oYz/lrFAtKr2Jx1xp5SnXnwVF5C3xq2mhmJygnnpeLPBq4Zp/eTp+K+S+mQpukBi8vn42VQauf/e
cxjMIne7UcChp8I3NK9Jgq5eeV/tMdn3MYqkhAFOGz8tuWlsIolFApxY5v/3Rrk3kxXbZh+m0qwy
7KVKc0nXoHFLvXQ8juuNFqQMhjee8Z1GeEuvG8c0YPWNxvxAQY12kNk3Mayu2TrdBUifKj7ZyjyQ
mSA36NK/LEHeMgwN0+7UkQY9S6S2qS69xvQjrHNtXyt4WNQjQBxxZiFA8Sjncpmn4Em+k/HkpbLx
2LAVmfZNu9oMMdEon6G/DAP6Mf4BXBZ4I9XxfmhjVCAWJBpU64CwxqsgLkDZeXydNPCVJ05mVtPI
5zNShx5pavNcY6yB0Hu80JJZrrsIep1PYdEkVqafRyL4VQl5hcvP+bQ60TbPPpJFuY65Zu7pMlo/
2WrGlFz0jAqmQazwqtHS4Mx8FLcz6dJbH4Fro/jMw4YOeS052Mk5Ay2k3ORVWuh2ulUCLahL89Ze
4UuXWe3zqsw7N7q24RP7gLDas2CZnextN5yY+vlCyw4B5tWQCBRrKauGG353eBJG3OAPkXx5gUl8
OuZ+E3wutdJIhiq7XpCUv7/pRpRBir9D6muExweAnykelhPyYpLjqHOT5wiJqZsdesKZFYr/CHHa
o6rLh+pUEdvRRLDX36v2PIpxO7V3Gsy//e5pXlMtI/wJie2IZ33FpRxlFC7Tf7+mcCC6KiOWYsbL
Ee0Ium+jH8uy4utBYu4AORvvKWIKCqn9HYWgaHc02EGHVDtbHHHYep7uotU70vZPfFN+OHis0yWy
D1A2CjDUCAykvcYVCITT2FJpO/SONIeT2Da3tVj70z+lSdOrBhcpAZn8P/J3NBkQ1ytp7S8wtxsW
n09rB+QEn9NB/WUYuqeF845oBdmaJqUWhTGLh5S6uXAZb2ioWzUsV1hvXXvp2CEgwU7MfGBA2IKj
UJ6oWDX/b/oAvRs5wpoR0GFLCn3xysrjXh7/5yn8boyBPCe0M0XAjbZ2Q/5uhk2vOCgYnHRb7ZYi
E+ob/fGJv78S+kwZwcEityT6u9KJoeoeLFNsTTFqGSChMuDLRVyLnDdYj9ndKP99165SpyM15ET8
sEKpsOsVX/asYu1M3okGvupL93eE0aJi702ujht5FMcV3Pfrs2CForU6MuWVETS00vQk+hEgO7fL
2bI2uSlLUQjg5MjneXcYBJb6i7QfbksIGHZP8UOm0x10phFZO0T1jj+aesc+Bftulm4fUqKDP3zE
1xCyLdZPNOCqAbLyGFCUg+4SEQ/KTCOUotpwLaY7hxCx5fnZZtq7Rn3awJxSvlscOVF3ZNah3dWA
T9WOplWz4VkqPx1X5DtWnLz0Y6yzkJ43ZZuKCjMwvMW9XxRfBLnpdC8f+oJFiO+2sHafjRpbq9xL
7Dkfer/cbMpQtBeghio98UcSR8sFJyjzMdWascYI1kxxpsufJMqlQJ6LxxmmPTHhTyFFYH022Mut
t+kRIm2E6t3bBwdaorgVGAmww6FprnJQysKMrGUDqLlq8fd1AD0gYUDhsb8MHLGpxMvUsfWP+vFP
BPSSCidc2lhhIR+2UV+B/+QAYQBbT1zau9GfSUvpigmrv8EeP6/e8BWsBrPIXevxPevfrSrj1Axi
T+np8xp65IHlKya15WhKUnta63yVBStSXmTcPYg4BDUv7v9cdoZOgPNvqjAbMV0vQ4rhpCtonmM0
a3LVNOHJGmdLJKgKuT2OOsw8H6ctBfWQf3LVzNUwv4xdv8lL32ko7UiI0/W/qidNfQn5mkZtd7fQ
pfrMX0e+TZjq/MTBJhA2Gd+MT3+jdSO63//CNRBr4/EJ8aJQUYEVdfnlv4dfo4bWMBOJDskmLDMr
5v2zJA8vubcN5wOiHb2toxSkFGeLlisGdukrO54avq5twr7Gyw37k4r+h6gI6EBPvtqoHm8twLTj
XmBkkZ/WP8xA0Yu+e/plo2qPjog0uLa17MQbPnuruS9vP1kB6NMfKPe1MLQpa7modZCptlLy3WQy
7vvciHxJ56N6G1egFj7GnASGPgxIveMX0pEzknl9YOwnyyxWxh9fYJG7VCh6E4YjYMM8NSDsBBPW
UGpB94rdjfopvRmxMk2Uf9tXheLR1t5wfA1pB5Gm99ox7dxMmYfmjjDw3hP50Ov+gZkU3hEhd1jl
Olrqxpq38xk7tOfIh8FE2TFN2ttXd1zhX+3wtEEAOBvDR3J0qnLhE8WCYKgkwdBC86WC/NSgfzr/
2UKLe04BewGstRsqOMJ9CeyV+rjDxLkiNFfjRN48QyUrD4IIShbgFUCnkg+qdK/3hj4D4XZqsoRU
0yqbkyOldoFlHdD7ajbAGnxxlNigwgDaLWNEVbSKc378ESot5WKUXCg2k4+jdqne6DgZqLlNdELx
CfXr2wdWLjFfodv/hR17HXDee40Q75Bp1buJoJ/taV/Pa1c5nqSUSf1REe7IdFmwiDqgbrbHwXTB
3t28D5WieOpIh/p/K7NNctSLVol3cFCSeOh2yfUwGYCZPxxvMDS2Q8cP4a31bB9fqE5nWxIHxGPW
nhH4kMXUZ304x2xR03DnhFmcMYWIgrT6fK4WtTGpXFxQ2NJF8TG0Yi94oq9WKpnYjhUefTmLWzM4
3tTYyo7+fUutNlJ/LhtfHbTIXXcNhbP2G0L2gSXOjmhNIChvl2dSYMCyaObx4AhMvM+qep+AIOq0
aoM5FVgNctlGS/avTordN8UPEFSuhSeJKTGeZ41wt1npYO8EQ+nJ0U4NAgqlpwJCGbx82YLqqC+c
F3scJeaKVIEOUFpU/2/09I0dS4SCiw+YZ6zGY9guAnVJniBBkp4X62W1KFDUcrkKVsSkWnvKaagy
1cY8KbcWsAbEYmWVcejuSJ7dLkVeDrCKG7bjyau5hiIJeH/cAdk7C+VDbf31ZK/Zqg/xKNEo5kBW
KWDd/6EyQadPUI40inVcthjkpYxUzxgcX4iQqGKjesMzgimnyt/M9qDj9WXEkxEzKtIr5JLxrbXe
+3M3Q0UtfcK9UV1QyplhnXbqpBn1iMQVkwo42/5nwS4UcTIyJeC9FJqHcv0gy2TrpfuUs0zVSxg8
ChRe+FNjZL7cfyOisAVoj+gkvdDyElsDs+t2hst2CYC/h3uVIMzg3w7j32gMHKJS8fEJdcRGOHNK
zHIU7FnO4TmWA7vtk8+IOuDMUqI8s3AXje9Q4HYnZk9FW/C8wQo9cp9zFu11pT23mfxiVmwQk+Bt
t/y8v9M5LbcVaCtdH+UdLkUXzkifZQoo2vNew9gZtHM0OunhWev4iEp7dVWTeGeZnvam0O1MifRr
7MeLuEXxreFC7f3G6Nhfk+OYjK6kP/BLKOI8dTz/7r9ONq8AgFv+B9AE15jGwBX2MBvB6xBw1Q6T
TzTnZp10ZM+jJ7r+y8n+r8l3ZBuPWtrFjDA9T+COPj7Z/CAkjQt3LMoq9VSUeBMgCkQ3HVm76/8J
0Zney+BIG3LxQsnSVZI19Jrrj5/WGusLa1lxMW3mrq8P5ya5r6zrNVYP7eVC9IyIviCCcWtHw/nE
ni8qsDAI7LY+D6pkfac8q9NAhQ6PlNp2r1Xd20iAawaQ7m6hcGZad+HbCxriFs86QzzDhHCdHrfb
doEIKBG9BwsCQiPbLUSStbuSate8jk98u1s6nDQdfFPVF63hI+wYcN6/cGTuJcVXAfyZ8kBPd9M7
JhadYujvZercIsNhrrJze9oQrXSYgnQZOLtsARMFlEfm75+zQ4P8vveX+FdRZX1l0EUhtUYUplh9
swnjBA+iKQqEKvIEDo6ESXIJG9eBen1vSXxs+rnMcm/vZmqaWLfgv9luUwi9p+Otb9M0Rtv+aWE9
cFcRowNKcZJ1/atQ1ndsbWcy401MoRKHQACl/RQJ4f9mPpFi6Kz2mJydxheps5oWGhMdAaYvWGrb
Br/qwQKxHttykol4f30UQK7JsOZ4G7pBefrrYt2CapnqBL4Jkj/OLv9g3ePEfUz6NYiBgorM2cox
2+vUIGEictfTmMhP6FxRI3DwNlOQ9cyCZKKNomk+gDiFqxHjBk3CDZyJNbq/jR45gATo1ycq9NAr
fhxJkDDputDies2UdE9NF3466hmsm9YykMqUD+EPo4jHks/o2VkXWfnp3ExNevLHtKwJ3gbGNoqX
IBa1Q9+SA11KSx95SzQnkmsudOCr6RQfkio5QnbTm/6Rmpta22f3OmDdDs3DFLHeU86RzUiVYGnS
Sde0XaLQfnTlly94rH9HmJ2Yo0Btv1g2ujF9Jai56a0Y0eLoWQVXw5WhHVDWDDi1AMg+vDuK2Rhi
TioVnGjRIM9XhlZolzu5aa2S10GQY8Oe1n6nLtcxPq6TNc2n7xqggyAPyKCMuz4RkD+57ANSngiS
p9L8MQk1troW2jEPSCzMZCCrI3z1UTHSMHOw1Sf+trI14uJkwUTLkDh/eFGiWbfnvu0rS9w8xX32
sqZslSNnxiYOb3vf8p2h+eUemcSMDag4vOKJP+dmpNfNRXuv0BurY6gN8MuAGIe5ClRLIbOyFQGx
bPf900eQEnA6aDHg0xd9v5Bej/QOxJgwYscCa9E3qXjX3JKcGEinoOhJh8bGi/a7M8B1qdHJxjdD
ChovuXBk63ha4FCH1GF/rnwJQpTW0+OTxkkK2gprshnqgiPQ7B5+Oej49S8Ch9qGrMZDiNseljDn
/ij4YTsoWiv0VVE54/olfDfN6EpAV6a6psHYVlBk9eT5Zvy+lXfVYa5pTgJZo3D1nvGWwlymAu/M
9D/PKOoDRQRVZNcmknEJev0v/jTOdMJ0zxINJJL9BXkQ/G3ygDfbmUv/vxNJzFNSaesx2PyEqdAd
XKkeh4HG0MtosyEv9zORKh/s6fo/JFTpG56MU22p148hRfgNj02QXDhnjG7T08/9RCinYUNDpNic
mC2qt7YLv0u3BVX2VS/DqQSzXEtkU8l4tDpc6AgI3uVnqPDtDMgPqmvM0hBO+ELCUiVWOHN50XXZ
cw3L9d0YvmM1zE/TbHbn3LNds1LD0n2ITe6amEWmuPfqaLp9GWKxW7ZkNTOZpsnn2y7DgF824fho
Zq44dJmR0/QkpmMWmq7qeDp42CfhnlhTiDdBzxzFy25dJ7atua11qALoWY+0tiM3dwe0qCsxb36C
21ETxhuMv7RKpJ6BB96Fizyqzr857QNJhPCpUsWjG4NXs0JpL5BYxQiqQXYDKbUXRORfqZd3ONRM
o7nBtKg8urMVKww6+XMy2lncMVd20hgAYblOIWXqdleFzdPA/WN+96aeFvXOhSlM4xa+kv/P8o+A
mYF9sAxxXBdHm2z/xdrsk6Pleueh3UO0gajr8OLQpURgE0ImN0Rl7bI/WDayD5uJyroibHnrFH0T
DAmsoecE2/MSKuc1+/sTA8QWeE4R4ONafDghtFm3YW/Au4ifEUFSLbufOQYydgdikclNJNeSuTf/
TV8YQrLPcMn7LPwmSXiiBAiMC+pf4z0CBai1SLgkwFE8raG8JrVaciXVGgknmxNT4wLLyRjOqTzt
U3eKDaJv4M2rtSniaBmqe0PtHpSnCmIQR7Swa8gtIJ4XD5pjNrnGKMwq95yTiePvg1nEjDQC0hqz
Y/AwgwlGlTGsOxr2MDPbtY8CZXvBdjWTA7FSTXel0Aw026ofJFPhNo77pIyy8+mLFSidy5fCS5ya
e1vLuaTrTHNZig0+HCVL4yYF4WGWqTpYFJ4RQ6ziwkje4T7zDEf6XbSUkmWFUvvFIJfoLQXXObwl
1fcX0vCqfl//44tm/gTM3vL4G6oF4d0O2GZhsLzIaBKPFFxOqVfp6LYrFncpRTOJeWcxluvbMxSo
m8UQvPiOz1Aet0dRCXPKtCgiplJj1csf5Wo+7Yn0bpWsveCD3iJAAJamSelRKzHb1/96v94WOJNy
UQ0IqTYBWaD0j98SRa7izeCN3rxIjLa0gdnXRvZyy8GF8mJmRYLtis7X/fU7gHAlXykL2nIMiq3d
XPe+mQCSMcV7O9qjMIfy1t8xg6o3Fvto9dmptLSNo6Hm6nrgMwpXFPvFTa7CPDjrzVLFGKdDFXJQ
dA0nUQ+3vdZwKlFyf/UA2TdpSE46sQ1wb5IrFvvAtrmLp2DadcGZvBfqz6gNTv4MKhlaoSBMu/aE
CdfL7p+S4tUu5EcCMuIKARzjFVRh0xyrGwK+9SW8FVTW+gH5Y2q4OTuzykghwK9L0InOnfuNe/jy
+4mf1sRzgxVopsyvvOGt1J+bY0Vg6ZHI+m0FkfpT+O/HAGOaZEIOdOpP1yp6rT0ksPCoMZF5SfxW
KtURGKo1ZVd3bc1ui4rfcx12mXhMsNZXBl74TP/HT8KHkpHVSM5qAySmkX6yqVhhQePrgiF1p+b+
mqUqozxjh+BmI7Bb0n1qmWQGq824Ms/uBNS8gUXb8MNf14YiClSnG8vlaflAvdEqJLGBPPtGeGle
x6UfO3qa57A8iO4rn9KwPUeEgj+nMSCHOdPKc3ZOSBpUh/GfG4iB0MkXFBuYxJUQ+dLe9GPjkn7L
GmGzafsbO6R537L2K8jr5A7ccKhwuzJ0DJ4RWlgcBl54/CQjr6FgxG4D7rALWttt0UVFT5/ijKgY
6/4RjdSdhbuNsui0QAnwdY355piwZfGSl2wT34XyMy4Gd+JgEkNqz5AZ/XvRFz/f+lJduhUtcGIf
PXVh1M9K9iJglL43C9sAibhClIpUWODhzTpAZvWk2TZqhIKhxEirLiMWpmtHjA+NfgrKwMhpHBAv
OybzXVBQf6GdTzgKJZ6obahAgXjrjn9uqtzHmVh2kVAe0/RLorIpYoTFCL6Bza9MG+8frCIXvcQm
tkbS8d3EQ3zAmQPGd3BOkWarD+xqzk1Ik+8P/sSuWRLxm01LP1i54G1gRSypCDjSpA5I3k1qBmE7
XiB+U/R0IsQbgU/JwiP5O3vIY1ZDp32jYlnGhx7/FpE1rWwO/shs9dayHsyd6D3e0Kdk9HfsrAVa
/aolAKd4T7f0VFBDfVzEgzNqi1Dh3SAG5m6nunY5C6vng2PbFG10PQKPD+rBQVxxy4pWMPdpImTf
RsEyVhYK5rO7Rv16xBFfy6nZBBmE48CqKOzhGhENAJ5aKALrROODss/9GxZrMF3GpjlIcF9tJWqX
uPHkP+UEEmM93KkjRD+HDWV8VpyWTEqjNSLIy4cYkyqqS7qtdzubag7viOEFEyAkGp5Q3iw77Fk1
rp7Rzg1gN6Mg9PXEW2YtdHBxrPPUB30kDcGzHFzY9OD+wUYQb0+Bt3ohE4CIt1O7IpDCNffW5nC9
v1BB8YqhmAiUXsgYhZlkBildLN+KPWnAodDdxweE2TSDD8XQScv5tP0JawxJggFB/6GvtDU8T5os
JM2jK8RQnuO18WrsJoDNOrczMcmHlxmXrq78fM2QGAwCO7sxwct/lJVKnAf4amY7+QsW3pb7HFpc
T91jnOn/b2Vkk0j6GvRIqQYFsUiLP2E7kdwd0owTpwx8wJ/rw/MU0uv3awNdgIuC1lkpIDqWAxsz
a6tJGGfgVDlhcqTWHEb4GHjHCc3fTIeL17oSe3qLOwsnq366zH3JEvmKBHwHQGKTo6saJ/MlPuWx
vKSwkxJb01DwTNTY5aeBaAxhQWXEpdQe0zEMZcyMySYYF9xFtjaNfGukw1AwxRxwoTqjLtlATDKi
tOP2rM41uT6FQcnA6mDzy8RoXjpYVjDrG7q6/+6OLA9BmVCBTCCjdOSCyiL3dhHb5oILyv/1mg//
gUEL03vHIMPIzKnvLMP1WhdL08KPIBGgOmGPnN9A2zNLW9527vCEbsm+TINRZqvCC1nv30+4QXZ2
qclil/BIfQ3j2loUTPeXxkIOYS0BF+PBK5YriJzzvomENRsoG6xpB18L+/6nZPs7VvGe0eddhQB3
cCD16P4OStONb5gpONYXkWjeC8ghrn1ptqq0o+hpBtmEiDNiqHcddkcowjg103EAHRObCVGlYPA1
w44Goai7Q/Z9xxBHKgOEf/6sYy73XOO2nqQ3WxebbSMehFWCQy2MK/EnR2spDdY9Y48GhObFFK+5
ZG3eP3ZohTwPwdIq5ua4AdRodk2gZA+kHUpJIhysOmVViBQmOy2Y0gXgylHU4r6d96gHpUTEtLW0
8c62T9UzvVz9g+IP5I/+0j2NRoZ3gZrgJ6Wi+VOhTVxuhGrAIUwMXdAmdU9FEDiUZzTncgY6+Hxp
/NpNZocdyzLD7gvFrQwt/tfhKned3JWdHDDq0R7+txKANfgVqOs8gL3ELNawMATwwrkWFLBlsbxI
Gx/n/8HUIyq5WZsOuS965qMlXPcyXQlKpyAciEywtCQfT4XdHAkTD41v4DBVAsop7FsfzOd8cI1t
0F6E5DZizRE02NdsLRPquG1pWoD084qhU7ZrwmTMdsrflc0Jtd2oIsGx6tqGDgJVQgfvXubwwnxP
HJ66rfMin9C80tOpOoAJdSiMNoc4B6IoXkKQYBy5wQxx0ysbLq3FQ1799trtD36T43mgk6YipAvf
FRgZwikfRtap++4a32fPI17u5+Qlustq0WWEUn8C8Ebn3EYOpKJn8hFz/5r1t3O7DKZFI7U8UUvP
0kYs6U4XdojCDROwnH+myc3Cvz2bzQsOl0HHC+1WR1omMzTP+oehwGjdCJlfCiKN8No2ouFMWw5k
OHW4Ba6Oa1qCF2jSfEWuKcTx9WxE1nY/CTfiCFIh5jr1+qCxwcZy1zW5P/TZvQACW4IYHw1H3zxq
tNL/HAYDzazohgIhwfXSS6JdXkIv9d0xltdqSy/2H5gaAlvqA1S7IScU9/vUrPPdaXWx/BU36Cc9
NxAoi/jecq0EERGrjSpRaDa/BbHKzjD+3fZyemHl+7+JA2BYpQZPnFV/5o4Do9baBHjpy8FWlAQV
I8SKIRJ3m4aw5Sn/Vf7cHtH01pFOHCCO6Td4G844d5TBeu21l2sj8U9UGfQsLuR4drqOjgUwvRLw
Cpcj2bPMwQ8iYOOFPRQKiUg9kqZu5pIvqYuBMEuerqRyz7mr9ELEVw6zUFoIsBxkejmT4lTL5KU9
VyG0XswXZfJjnqDWYltCyPvbDss4dcTC/stuhjKrVoWs2g1FvYohsirQ35ToLWnLuuDAlyU7sQw+
OEvAuNkh/zRShkieKRlzjPFIjbjJR1yMPk1AcmJDjIpDfzhC4XiMQeebgL310NDYm7EF4+pYlY9F
vALp/wvAcPP9CyGiaRXI9OJvgJaL4fN66xNKue66x93wKJ+DMm9o+TF4+/bhSkaQnaZ02hzaj1iG
DeozO0Pt7K1n3woVTOUanPe6ZIe9RTBeldOloAL4XIBb0NVwez7jh4VvEEfhCC0gOTQsqe07eROm
uOtgBFcnGw8/ieVow622yAqUbv/W7QNtCJ4iW03h39N0jjwc+/oqne72CdZ5VgD1L521N74kitou
M8VXGB7GbM2/h8/p1166SHz6sufzB9cTMTk+5eEijFAsN0wsvJ5MAQ6KXGqwOhZOX8Oua0v1Ngny
jaJPFSpoSUXlAd8zPUKyqr5QdS9qvX5gnpGMFqDPvUFH4dHY1wG9RsD3Bv9uYC+SZVYH+3HS5CRx
psQ7jxoqFgO8zAZ+w7n9Ypn0ZAalydnAQ0uSWe9eucJDwHiyRZBj9taGF9sdpdzPNa/GRaDk94JM
a8RrMgCxJhDURTQE9iMX040pDoQ04iIznpS8yl3y9mAPpskp/HiiWZLTMLxad1P+ouAMeIrVMgS9
JJi87Kdya3U6LzoCYhnNq/oGcoVfIslghku8gzMW2PyM5Ptuf8da6vl8U36sv41wlrOZlm9SXMoa
5BG9aBVONtVMppDGfH7JQDvnyvzS9VITfTQsiYKnyMRSwcKj/V8ZZlObHiv6sJNe4QqHWmGnhQxL
OsAtELYcgzqD1Eizl3pEmlNA7gDW1lEpHBCSfacBSjRpvAOC0I3RIlFdWY7B8Y43Ab3kpnCmfrg8
m136BzBSIQucSR/9B2UOvlrf8kEyTUvHWTlYQJ0FskttuDXkK6XrIWpnA5MrfCXmxKG6sdcVyYOS
5Rw/rNyBWXrqWiSoSWZzTSLfIOupgH83cRnF76WNXKEL6tTs6TbTSTJ8Fk2cWfJ+N6gjtkdAMijV
cjYNeDh2o1DjV3CtzLbIqoI8Jhsfxwvstyok9pxHWOIgkqn6qvRw0FVqpw/l4FlgBCUk48D7NBqs
zI0QnGm5Kl6p9WXc8uCzXAtzJRu7m/TsGbGTpw198D7+6LPQAlf6q2ANFflti6c3a7Lm+tbxQTN9
ba29sj6wbJ1p2P1faFTzoAGMc7l/6hoXFrvWSBvgUxLeD5oUfhgYZSoW1qMyopVSgQOZjrVDTnbU
4RNmmxAvkTi9o33l802UFLd5dT5AsE5KR8ORmRjLmDJe7AYfFresUra9tgiRronmbahymXyQwbR+
vuWOV31egL1e9ye1C0uNhtQlFyvw4416pCebwUSGwdc0znZP/fIWe5GgNchTpsBQqCr7SqGmKtlI
kFpJm4MBgGL/DEeBZU2ccZcoRD4y8ID3I99ix6PyFS6mHV9fTp0QJYauJ8atKoSePW0dzS5Z4zZC
DZSRPZUo00Gx5myBGDv0OxgiQKEQs4Jg67RCpU8r+6Er+TMMJY7OUEbcpAkFcnGnMNr/XvB0UoC6
Kqn29fyE8piDCouL300ljV+vGUVPrgmEFNRrKLgTLg0bKm25oE5R8adEIMLjwXB7CB5KjGJEqXzb
mS1hm4UKWk/U6ijHezgjVcAOaS7RcPdWSOVxiQdPtpIAwHSdTUlqT3vB9hy4QyVfenVm90I7c11A
/A+4C6hoxuHqZd93L0HIa+X4hDhqY13xIIErRneGgtt6pBNGJllpc/HMPc5RuIres4R8JJC6tkTj
xFFAruePgeLlIEO24muUZSRRyUB182zpXJ7Q5hGUReC2Q6azsc40L/e9EzDGw8sFVeNIEyYdvPlf
KlyeaoGiPymW2r7TSTvY3zvgwfPsykOPxTLbzHYMoU3VeRqxjU+KGQIOBeuZfJdWxNqFe5/44VPV
z/RLnHDEwCsn2IM2bS8fbVYpAT++OWdeMrGNsBc4FTXtUuHxJ6sQ+dCVh2dB+/lyEzlJ5myxxAYk
Y0BcDfzaio84SPC8HS5hBAogpwemFWNDPzwipAG0h/tyCAYScSJzgZIBUIE7LsULk5dAbJq5s5zD
4CAwz/YD410ZTjjz419IJEequYho107zMK+z6u2oOOjW26cMTfHRMbkMNe7RvX8R9Efld4x4P85k
Rh1tULpR9EByMGIAKoOfp/nHIowlm7frHfYyhHEDJK3Fl2fmPxY7yNTBR7xOOxwj3kKQjgi9gQAd
rNCtAgEUhXMdXb420lxHThOuveudkai9mb2ksi9BJ1MRX+V9YQHY3R7Vf3aEV4hY0Q+4xRfuMkhh
MWp86a3NKcYVxLOp31e+4PJ7OqGdUY4akaxikuDhuhBwIQ6sJxlV1gm3jWWlwO9pOT9XhyyY0FaO
1kE5zUZiRQJ5C3cjXf7M7hJ1GLKxnFnQgJDMBOvT+rMdf9n4ta00G5zRGtsfm+4fx/D1PGMWO+2m
tlTnhF8eMWWKZesC5+kr/cueJq21JxeIVTiTomWeyaJyi0JBYxeEgs2wOBh2y6qa3MjhawxlUcbY
uLtqsF4xNiXBZioNvWFSpVJsFXXnuFjsGoBAHHA2tXc60J1bvY2mPeGf6MgbHgZ7EFMkjzMYA87w
tnIhSKzaal00kHO206yvt3UNkGGjF79f4+YW0TkmuZJP0QNp7eMSD14a/3jxCWLwk42Moc10S1Ig
Ej4qow5yluLzqqaBpoXJ5gDPerqWpy4DlrvfaVqJEsL8Sb3f0iV5ZC7miN1umaWzV25lmrrpxjn8
mQeDNggiH8am7eqI2+kq8lHHx8DpWgssM+qG9X8T5pNu+GJwm0pBdMNDB6ECEgQwxEAnexEv4JO8
008tFONM7yzpdrjlXZUlthCXRUUVryIVcLLndnkKJh2d0nPM+T0j7iDsHq/sHHRrTycJ0dvwW2RK
+jNdQag93A9ezCkY3mctusY+LsAi43pxtnW/fLnjh1A38Msyy2E9x8o29YGkM/HbhEdUs6MHlU4/
1DeBuzG5fDPhuygcdlNM5PQ4Y6iomJirojd2q5EnuPCBo48QHoQtBw8rOVdCHtZ/R0uWCaBGEOhB
JSSXtmWcLFWJ1xKVjKotvQInZ3pFekFoY7coeSEyscup8oZHmQwgIE3H9z9RDsQBgZri6dgZQX+W
Kw/HzjzomSyU6k7iNIAwe47IrJlxeoQo9bEypbEHGymdt2cAShj7jIqk0F8IVnRqBkVYqYElmIK0
VPKLZR19mnd4OXhtQg7y7HpW3N7tiiRbmE0yI6flY/fI6nrEHxS5VzwW7rVtnN5j0GgFeXqDrHhD
k+4gnAcoPW37yoqHx95lmJ91r4RcDmsSWtnqcZHMAscRE79HmRMFY5/XBmawLHVuYsppP2aVGkuB
/ZEaqsLTGwJdTN6x82w3rAcSogjuaoULweLYbMqTgaI42Ot8UYGCASP3h8RqZ/sqTAwqsZ/dIXpS
/xaON4mVJFnEAzE+Jqv0mT9CwHx7oguQVGGrL2Lm4i9ot+WZHjw+f27YTK6d00rx03tiVC6Lor/Y
DDgXvTSpqSJSx85VXBPpnkUYEFvOTnHWd6IANY/H2HoEKWuiZK0GvqRa+HwRgJPOuMs5GLB6LgsG
VhCJjBtxqcmn/9hdaiD2filzWP7J6HbPvCloHPaUC9uFoRc+sWtr5GuyW2MQMGeS7x7yN3KC2gt+
Ols3QpwYizEqE08hMwA4CzJnjvRZ7PYZNu9YbWm0aiIaVpAraNszNF0teG8raYdssK1sz3lIzUCu
JtKAdaL6X1G+pSy5XwUo2KNJCcUbDA+BT70K96IrlbqVl1u5Fubqo6B7noUGjG8dveLo8+uf9szD
97n6dPNiIMLX6aXXu5iFBJ9J0Rncgnij/PMlEzmlSqMcxGR5Ho1yvaZgdV1La4Rq+TVcn/hstCgS
nPLo0kstRQygjSU7S7IQJRi+VrcU6bQzdWST/fRItpkpKOKNVQEFt46r3IF/8XJUwRBWW5VY6nVc
ken8c/SqrtzKStl1h/L05UV4fp9s0tFVOKEUR1AZ8hIMhML54QKZiKWZNAawsb6LceVPrzjocVYY
31wkFHPvAXDmkAbQ4KgtKrw6xZ9QZNbYAApyC60pjo7pNrk5LInhUpdhrXWMlpf0RrRSz9k3482e
YmD6QCWzNgSgflQ54ZjHMGOLxWhlVCOFTbM2Kz3G7CLqzxmWXtdizCIMrNP79b0rhCsj24cBXju6
v/GMikCtwTH2/yfj2N3/jXzTwj0tE7HwkMYy5/vft/mMzwx0ktjj39+EGcjQbhRtcRlNWGot0N1h
STGfU3slBfxbJog3t6AAHLb7ry6AbnWOLS3CrhM3DE4zWpi1Z9KcMOk+3hYoy+gJdjpqjavMww+J
GTG55z5TOgkK++2Jf8/4+sPuM8WA7fKviebpIO7LNAF2XIglhcSHfl9ihpmTd0gNf4+ATH3p+E8y
JsQHZdUW+w1hVik7OOZC+9VobNTRnlaOEJfjcSuRueODiHLkUkzAofkWxiBSKRagyjNq/FVnOqgd
cuITkslQ5V1GP+6bOHelI8ZeC5fgr8unTxAN7CCkZKQgXZCA+hd6Nwggd8SawEuH7GW0sKU5haYu
h7BAIII7Z1mxV3Ps1JirY1kfFJ98HKlxmv+j1MB810st/4DeByc+4wRHlwMwi5/ZeuMZgxep8Wxw
uP09bAqOIfNFyzwTA3TMmgcl+1MpoZOIA+8ejPUnFmWxQpLqnJyX0WXNxHX7NzvwYKpWI65LMev0
wU1EjLqjgrRnFnNaNcxh0oyFOc/tS6VpA4fANhXxsG5mQ5SCIkT87nttYSseQWGcxuDkoZGlAJRv
Lv/a4EPUqAVDda64IeSARQUExZtmnNiUus34lL4+6vQJjgNS7AlmIJuaALcjW3A+h6LctS+1CzVe
uFswhWchY0JnCS7Tq/+OBQFc7FZRqhg6aHMMPIyMRdMT0S4VSC8d/AhRYTlL6ZNfvgc75QFeFDvW
+SSMhCkuBC1TiqXDGhBBXfnu/emr+H9GLobRUuRHUbSbo3CWyKnU+K4oxWHro0ARadAJRkudvNl0
Vh10YmD0neNWk1EBTDZv430fYRADAXaN2maFOZUG8JwM5brl8zDx7LcpzQyAbz7mwJ2HQN6OiDnW
oPkj0Fn7KXuQBDynNERlQp2pJuCfYZlruK56RV9riqnGtUKf18BWj5luYfOa6JQVBnDbJM45UBx8
JT/MSeposaC5sxN6txtLzOpf5M+zAOFaCO2YDzECnbs3vD0fTZooQqvh/cmomoCIxphzIFtGdIM5
ah/1i+j5omBRLIYOrZN1liiDl2Pt+gWarEHt/PS2kv7Pnh2edyWT/4wNq3qWKRDEdnmm4SHEcsyA
w4lyjhK//xNaum//ISCKwaIC4FTWRmLTpqtl1ao8539NE7DfUG0rjwNur/4hmEekH+KzRTVusqVU
VksgYh9bj5EaHpKipIZ6CT/Tq8+SyXcUv4qo0DKQjgy8AAHDzSqpnaz8/G3t71ZiLQDvnV+GBp5Z
RVMfRAr6nOI8MauccSNCaArViuHxCsVhWmYuuhdOzCW4fM967zsOyCK+QW2JtQjpmsJys26T8cje
vk4xjtSJO/onOo3WcIz5Q+yEQIGGkkeIHxEwkeRzo1HzV6598H0Mat58q1AQb4i06ZZxercAb86p
+x/sn4eQl4Kg3LtioYhgtGsCO/zBPzJ9hKPZCBCTnUoR+DbJZ1HIWDf0w7z6bZqs0tLcsmmAJlgz
TFW6UkJUMnRqhJPIu06g+zHGexdC1rvvA7/vbnRfGB5/c8zVX7R9UbC9RKLTj375LWRHYptWleW1
FolR3eyd+3HIb6Ru4a3pI/gql0t7x2tTZEyVASrMjv7c30xNfxTVhYvsPEEObu2bNtJFwMRwE9Z6
6IGqmk478uidKqNjRVMlOK2tBXyeDNQrZIoauwL/kygD8U2zkOVxT74Pi+eZok4G1/UosJqYC4h0
dNpJf+zTvydR8lbAeRo6BxaAEKoEDhYiD8TArEep+5HRecMmrW5w06r3DjW+6Vz0QgptKOW6ibCY
g236TwEGqNe/mFbH3f9N6JVQKRp9uqN9rgiDi4BvcsokmmJ6HXTaK0+VYs8oGkLm9jM1wQIqXlCj
MDo76gugT8C446SVj/dTfrKt1JIJpjrc/GzeZ/46OaLN+Ci0lnJa2qaf5EavVPvsCnl3giQqf5w5
gKAhrzdpiHSFwddxXMvz8uO9KedXXWCAILBnqQYqkBt+RBUEinUHmK9iGC4Bt0iCb2R0H/gHX8Tn
3DGCFoh6bNNHYRUSzp3mzMFM3rA7hoBeU/oOa/WApI/wJsnhH8SgCnCEqzJClnrtmkVDjyIqdiiT
s1F0JdNfe3FY7zeObp5KHSuSZKgXToo0KLr+MdeRQ8XDYzNJTjrQa885r7zw6sdIa8Ia0VJzgS17
RFOPHTesUAPyJeycBhE59GAijLzxj4Upw49RLsGKoc7nzBUIB9S+yRl+3e5nZKNBsJ91BltM0ucB
h2puPYKOxvNBvM4uIgiFrS17SfCc/fHPY1N6EUmefhfRLcm1AjUbPHt98awhwxwrGZykJGKZASPA
b/8P4y8R0YyW96UFTQGIwFmQ+ZcnSaYghjpL0BPXcPG7gaAUfwmL2VX1il+wex9kvXtqqvtfkCFt
dYpxcItoGkS5T2ZwOYgiRYk1N2uiN4FQKbc2jZAtLgk5+kcylLznTd1SXTtcj9szXatKMTBEPRdU
aZmpkUMiYNQIrnLKMAH9/uYbgfF7AdBtyjf4fvxgGIrM+WLIDWAMd2D5iLEZCNGoWrlqBe/viTv3
ca8anHidyb/ZoZMBZe6FqbLUBOOabGydcRzC2dvE+yYky2KcjWvtlPVDgi2ZhwcHovpU2OK51oHe
vlDuSWoSbFwl9YRCB7uJYtRAKRJWtsbfCtzbn2w1esIWhne9mfRya+FIlP8omg0X727hIgOGEjXD
YIZiLI/QyQ+z723ahbHaBjRwbSy41692lXv2mrmn0VQ2GRFojqhd9HhqFOBgxPNwo3NFg0vch9Q8
b9ifF0c/yZv5rjgaYkf+x2JpRqIu1ZRDkqMs/r8IApQINY75royrKz0Bdf2OYZuwUk8VQXlO1N13
i8KAfn+EJGQz9Qy3w44yoVh721TJ+a7ggDYLmuvrGDKBuF+lqBSNrfefGb5WOPRO7I4N9TQieQdy
jLrLX5VaXCI2+UkkyYLjprnmPvFlXABmhCkPTwnR0Jaqcb9kDoWjCZWz2qT/6BQrYxiV5ANyD5KE
Cr4NveKJUOzRRY9y+gpDU1Ff5DWKO1ak6bfVtp4cJDlM/po8eCMnXA32VoLu/ew+k7Wveiq4rLVV
ljzaciuDopt2glj9KeNuosTznOyLPsz+hri8gWeR0tmV37+gqcka8uYjB+KaLgqStGX/S2I0/vDT
PmG4a/FE6bbD7uaWAkhk1z6X1WLXKKYmjn0OILln3LThc/UGNUr77BE4i6ZZxxtbMYxFkawe1Pqq
VqKugd21JN92x5sxbiSkRzQQQTnbR3h3YlqICzCV2H2uLlfjfd5URZwNGUuPP8Q4JR24s8Wc9Q04
spkzxtA3mWKTaXEGr81Fde8miKDI91HADLQFMutMfIHDVgZTRmQhTvsRbfq5TM85LxZ1ozGyD7Q3
1hdDgYYrxn8BzVZUem3Svtfy+3iJ8U8zBF1QyiDSFwyjbtWLA8GCx/r9PeGLMwAjCQFrOdhyp0Xx
rkz+9gXLVF/KTP0N8dlnQ89uQnqtrLcLxATGytvTbvxfxECWC1/rggvby8BCNH2Wyiww0oaJAtTB
+mWd7eKRxSvwzcLUYMxT0eyne1g8wl/GDusRomys8QgWUJhTW3pIA1MQkAjI2k9ggBlschdtfPf1
+g+YMAB/mibYGPdFxyM2t5+USjFQjNbLca7gHNXNo9xPZaBn9TFX04AjymzCHExMCLgxwS+m5WSP
FMhuR0eeDmkOdbhk3cyBphZm0Fw30fU+rQTvyM9oRq2NdEBsvNJ+Ijq8weW0DXA7q52JKxjEQ9SF
6kLAtb2TAkrhxv+xDZVwrqMDrg60MzTiLTjk1ItWGzwQKG2A/QRlAygcjV+sUCXMF2RXLI1YnAf8
Ke2FPUJAaMiqqEGyakl1DVe2ROZP024wfWTm7tD8qVlrHAbYldXDAi3W5meLzHmcuXRnuv2OdApw
o3LIiGI9SKPhs/LSUpWGUE1Dm1YYYDRaV2drr4dR4XVrCZHPpYO4mon33dmMcd93IHWQSCXL9B/L
4nWusGrIlDpygw6TnuV2gcwnob7Pvto1uuJ4h5+WOXRpnWRb6p2490nt7rAjSnRnKGBse3jvBT8r
m9UTZ7vIaWmC8X0ptAFZLa30jHV1teprcOuXe/oiOREAdWrK1OUnr/2UMFVgk03otBVr3ylB3xID
hB7CCiYRnjxGq1WIJjmicK20SPXMrC+wZQo6QR2Q4LiP8wZc8RZoLM+KSUkoVW9TygHEKlc0UWHx
WruJyKS/U2hZmN0uYGKtPgbRKrjmFsxiyT58aOcoIEFwBcrV0Q/sTRPqoVkoiQU+VBgebgF6xXmF
K2MNPmHrZNKnNV3GAOJIkPVfSdc7MuTk+xbRHMkT4asoQxEXqzHwkNJHUficNmue7RM+dgxrKnDO
g69P+Ybk35keLjIvxqRbCT3THpjqE+k47kHZudZ61ep4MaSX1PI4cHInrQ1z1UMzsgBoXVr+aXXy
psK7/7nCgVbn5uS4FtprQH+TZWhNDRqw1Wk7p8k9F3VLv+Vdj7xjtRIbW6RjrObZrGLnk+9FWMqN
Co6JXgUgU58cDtd4agLC7yqjOvpvkUKIbCfoTY1bfQ9G3FABRGJBmY24nhXV5kpb8FTHNIZ/zmdi
fBv7lDzol66LOPEmSQ4sgaJGjhUzzxXTlJDlgrSL7LbQr8b8D13l+UYr+EV4FFS4u65vOoBLMKfM
1xQnul4RhPpnDVactPvXC+e692117DS++AUoY1QgD6RDVY+BPEZlGuuGKhRA5ycWv1aXiO2sZAtA
Ep+1uhlFBCjsO5VhjbI7SeE5z3KDDjCPcpTQnYLatXoyJHRTeIbU3kFSNuqpSC8gDFQVMdqCVmzS
i+kayAhbNxioaYiRBgYaKe4VcWf3fJGifkxRwSlBrtjRz6hXiXWxka+D4wQfpLx1t074fAFRXBBx
dGVbcI56fEHWjaKxmmOqhBTzxdZczantkxONr/+MGVFVvhUK9m0oM24flPulfIvLFzKlVDqtlT7X
o+61h8z3dqKIw5FSDeK6ws2GlPKnYvb+d/O2nlFzKKeD03I1yoKj7BhTZ8wiCcCumbj33Oa63Tao
WjquYDoZ/tuptJXZrNj4yrpOGSny65LVK/gKB2DTJQqFUBzFM3jwfeNHgjf6V/JxSZUu5pro4jNN
sPGkty9EQtdpJW3cE0/Ct1aWR/+1+D00BtGJadQRYOVj6QbxLO57d6U3r8QuVr2WPJJxMICyEpp/
HRpE72F4nCrMcng4ry9Bk+7P/bgUYpY/f1TqjuEXFFMlR4R7Zjzei8busnNBQ6WmToMlZXerTlbf
ycs5Yiismtn5BZT8siaSV7UX8xphd539oJb1GxG0nVWdg8Lnf2KYJ/lSc3r65ODEd2+U4gLyu76M
ElKaRYisFHbTEGQ0fAruciehwdKt1krBxSjPgAvCcq+bxvsqqjb9VLzGDfExTOd5EqNRP8w3BUL4
TTZmr7Vgnf1ng4HSu+Cle/pEjONdcTCkUInna5qGGur5fN/ewzy5os0lGGS5/H3N35Q1Tl0wqRDU
E/iFWHtue4Ci6Iu+XWpZW1I1t5VOPJYhBpxzqF46wuFAoRB/SIJw65Jvkh1Rphpc5JkbYud2dK4J
IB9cmQnbzJ/ZyAKyDmueS9LOWBg6IqkzV2u4xnroBAtG0U64R6NFr7pnfZQ/P/seCQNulYp4dXhl
n2EX2j7ZX4MlTT8buOj3k5cUUVHMh4pK9bMaiSOZzs+Xj5ZQUGMoIaUG4EUDW0ifhWiKSmw21nhd
XYG9gDZyYEH9rldUTB1cMjH4M/5Vg086suFYTsqazJ7Yfd67vtRbr97xkvH4uAKZD+InkYybotvg
Tti7pCCN6r2Ek3M+iP19G8bYQ7sqtyQSdc/Ki+b6yR+SglxeNeFI28P054gzckIHG18LqPUaayFt
lkiNUCB1gkdnyq8kPmxE3vmL+YgkxSGtVTWa/ywGEbHTbYoK1L3aoHNFchqAENi/5vUf62M3+J7t
ircV8CphxHZ/7FUqMfVMo63T3x3ToN29PCoZZaCMml03y6UHlFO4r+8q+2Mbl1d8tj0bzy4ZP6KR
AXFFLYXTHlD2wQ1k0HTz5xB2pcdVVJ/9qN3tPn5mffGtxHJGHHDk08y+wAB4Uyl5wL3hT+bWSyR7
0eQj5+vCzRjekW1jDcest94rroAuI5dh0Zdtm2aWvblTnjDqzPV4JENqqggDI32zU3V4F9cR4ufR
vRhWQ1+98xWD4FERLM3TxWEHH3McrsawCYv77e5cb1u2000nkjudZnp2oaeVyOSHGW0rAq7twj2I
xNwl+mrZVqRghMkMiROdoVNqULly++GXl2omPIbPh7o17Yc7mHfKvJkYfpAPaoLtZEucl8GaOiId
MVwbAb4VL69+i0P9yEASqbl8GMdZuCAOdCFOTBZfVDJczTAO08j2Wv61nlSx4gjF0kqrJorBZ7rc
FEb7oy/ElBc8l11qkvL1aTTO14Gupk0IsFCk/Weo8C6Xao/QshtUcCpEkjZDr79Gq5CtjbxmBHY3
+qEigUZ45nsxUYsT66JCz1vv5dvqtiwzyPR/IJBnPtweuoAKdMQ9CXIyqvrBShi/P5v44du5+UVy
D0chDyS5F4eKIKFMN+XPiWQxqMNxXMD3rwvaNQSAN40SlBgaMObigAteKzW6zi3BYNDHpl+zr3kY
TvB9VZJ6tEcjkVmgHAA5m33ATzeE1IHCerZE9SsZsQWYQcf2CxUFkXEgGOqCQAyWO2mIP+Kcl6J/
mSLFa4SKIoMgVPKjz9a4MgJwxh3bdr/m721lUNrEUSYE0iO2gTJ5vJAOjNynCmhi1FUF3VdCKe3H
oHukK+jzjr8JDtfLQFOlJjDag8yCF62vJRUXsgZN2y6tSLWAjl0Y7RbGUb4yTvbI+UAN5ISJQrac
RJH4p/Sbs/08vexp5Yg+0Z7pdL2ruuE0zDCo8IKNEHLVuqFc+cmFqkF3md/ooFlF+gBjWpZZU5pH
8ObPWoN7jUacLsvU0aNahaudkjhsFryoCRm0NowQJ9/lK0euViwt4tlKPhtlQs9oFgiGf6Ow3TbJ
Eea/5MW1M3ODt+jusgex4crOKnoehyDapQTYbnWeiB7ixRX3vVF5tiCQAtNZEkwW6dIyF93uJH31
TI13pGbguD6rFAQtaFAkY6N15sgvkks3OzsX8qx933uN8KapTuqBjHRnq8lipe2LzaW5m/Af3+P3
rRGxoeNGPLIytEc1NSklVoBiop79yj87Xc5Sy5qj7dE7at+OYB6UTQi3LE/MavxG86tlMoFLErOy
ygYzkFlVmWaVCbjJmFQpBP71ILelhVkYrqVGetADyUEabGoWdKecdqFGgfhVY3i9iu/ZxxKNAK9h
RJDrjG1a6KEhcBRlhdwMQ6L5D6cBC8hzIs+9+0uqxag1nJCGhNVUAb0cx3Aef6OnIvVqk/OhgAnb
smG//HorxLDDbeOi0YiKwL43OaOYn9nSBUPd6zWQP6vDAHJeurSxbNn9/n1q3TQYHpPr4qwdr5Xz
bmrzVOczRuRVW+jUF0kWCv9tm+39w1Hr6Sq3oKCqzPuIv6W9eEcnuOx900DommrpEXgjFwhoqlt9
eT/BRAG4dNNuZVfg9iPCC5oEEwr9QYJlEjcpYvhq3CDQjrkZGboYwI9bvt8KqQRMcWKsyjQwq+Hf
v4EFS2VN9cAE8YhU7ofwRjJA0Cad22m4lfSop7yiIzLO5CXARImMInAHtLBET8PdgKxh52igdcXd
UM7wWAHRz7gMCHhdcOTZaFYSDUmdJYrhr7EHcomz/Lk/5RvzIwjmgJ7cabIvik8igs44f5SVBzCH
Kn/35VzrP83Ie03GJk74MDwWfkAK94Nx7dBh6akTXOcIG7NU4JaSR6/j+ECYdAwWB6M7Y1Cd+TNe
nET0UHN1mJlVQg5MhtQrzZEDrpyqfJT4RcIA4yAu40epewf9XWEirxC9bTWHy5xvbOJyDHSLOPs8
gAZhI2repLCpvYRkPdqBGXo5MLhAyl02z4z3rSU0gquIGR8d/BWogBisV9gWQTS4HPvbJpW88mVj
VvHEZykkwfYQsYEdlyNY1x+0YdndU1JQj57k1Ggq/gLkoWVlZAIuz5BB8bhw9uixsPYn4QWCslyG
jtFy1SICxgMqxoZWN51EC1y6O4qvnwFWUKvDRRhEWXPA4MI7mY+6OnMm5UlxEO/VMHujXHczib0H
iHxJUHVFZO0BmUNjor7Q0Egrb8sUsCtaC59tgpnEFLRMfimMvoVNpjVsIIZNnge/P2Ct91E79IMD
pDrzmSmLVd/0K9PzQjSsHGYOIvNR9AdAZVA9SbeD1QvEMaZYQ5Yhk71ht3Jb9weaEbFPnujmBGYr
t/BtOxxnRXX1xjHV1c5GwRTHj937iCDrppcXqozDdjK4dCjbKP/ihDDQaHviGn/hACbdL3kYDOTp
GxCFnUwl36WllDuec1xt3GLqKvH1b05Uu5PfYzRdbGLihwESMp/j3jf8GhN/n0kbbmM36+LpD17b
nU4TQCidh7ueHsDgWZwlHT9c2l4b2DROCcScIDSPFO1FB+Z7LQGjVEIkjZXQL3OA2c2trNR/uC/B
Es0QRsiAXF6KnOBmoTmz7XPNFB6hPAK1T6IMS95iC2E5Y+O+BDL5xgF5ccEy90YwfmNvkeTFTPFX
23//N6/bDQjvC7RQxjpYLUH575bF/oeY/bub/P3VONmV2bT9Ni4DanPVhhURMPPAD37y3maES0py
rBTbAQr+7z6ZUNrHBOT9SjEMqTzyHAPxg/UZ7HBiml9cDXWQ1yoSfQzRg/6MEKTOqDhfxIXyL93V
fgnio8rZJ21UoaXHVopj4Y+Fu2a3TbfKNYlNMRq44AEYFQrGWnblrKPkPseSnWZmTFQliVvvsYsD
gC8+VgP0iH/WrEi/68OICmIR/jZlfSRsTt850vfDHVtch7kQ+m2Gx5k6ri27S0hnv1hYPJW+KQLK
efmPWVhkZYwCCTO1tC362A3cPIAvXQazYzmKfs/Fk88nK5IyBL/m5pcyAJKI5/xx6jo3nh/Yqjjn
5HlsyveFJxDUnvllNnjHzXKlh4NJCYIOsRw+HAXP+Jo2YcPY5Y5EmVBvSgci2JwaqmuiF+RbXyeD
JjlLDkfFFbEpta8RHZk2msCWky5SFZkSijzgt777WJlolxdi3/wsNPtEKx7bqqMyg1/EvE/ezx3N
JQGO57rNcbF4GGhq9DrkXJcFaSIx/ndfc/nDitMeeJl3zftnUgCvStkHFETFq2hZcwXLSVTiVCb7
ce/ddrq+mbPFX2smjrpDVCgAZsMtb1iABnsr3gyh/RTh8VAKn5zAp+2oWE969IsTN3NmpU1yYr4V
ljecSrwHNXbaEdC222sVTswmhKjMlqdlB3eenoR0TN58HFqrAqk/OV5xYOfW7eaKchgQ3jfpPB5+
v0l3XEhZQ87a2DITKhQ0by9gZ8flbfQXWcHd9gIBj0X5494UcozIovDuZx7fzxIGL5es09E88Wqd
yh+cuR9FLMRlW6tUyUFdH/or645PFQqA/kgQ1FE3C5xf4c9vA/rrKQ8qgewhwYEFKQlr9lvIP94n
CG91mDBWHLunIX5APi2144QQunZefknf4bZFtOIOmUZ96iO/gG+CWYXjbU8U2ibv4qOPuOPyAzr4
JtgGfSAuo3mG8clHZXwyUvq+Ka0uMDja13De3Dy1zdAQOkL1A8y3gLKPqkyK7ovDgw9xyTgOuzWC
TQXt8+ylrB+3L8PjP3RpUm6roCUuPJg9+MFLppMNA9gtAVlYHoh27NlAWj/VbAsd+7oJsfUlJSMb
6xsDK3ttZXhrDlASB9JYZ+2vogxU73gbr58+M3lhUTl7orSeFmMslGTVQSvGDZyAgS68LSXv9tl3
YrBuR4qywOazJ91cgPQY63LIGP0UNkDUtYA4oUZzlPv9qVWlGGFLuUtRuoeL0nZAmvLKXOZHZqLq
3ADFjbcyISOV3cofdVBFa8VnYWxa63Y+B8kXi8nQOEC1+/OicMNIXpNaSTqTfNGAQYVqYoPQdxjk
dJB418Jh+XzoOWJoFBfiz+I3Ju8OP8ctvO9yItM6jBNdUTqzyLyh1aDbtz7XlDfw9HhEtwO/raJh
Yix7DzDwU9aBuomXu292lZpPsRAIVivFhsSevAp/7PwxdEDMIqKBTMn8IbDoxxOZgX6BWrhjsgf6
0IjZlnOzO1IYG5q1nHAql+zB3pLD13WnIKtN4fK5QWnrpRm5spM+kFQFth1t70A5ktfTvPk2P50H
Xp5q6S/YVVi2jNVd+52wtiYb869ZYySl+XDcG/nrXQEEpF0qZtMjRBUt+k3+dIcBAjtTSMqrFbRJ
nOwVmVPH7EnqXWbs5NL2ieXSNHMU+j3QLfYuVGXFywU+90uIZTQRysKoFdIDEtO6l2TglWIZqIry
QirRfHYmFyB3+AzTK7gvcMyYedZfUFCSNyd/gQuTc7rFTKeNSHw3ijbF171UhBJREk+zMxrLnf3m
krYD1yU5uA+iiU9CWqSQX3o3EQNuGADJ8YUgUDpQDuNkvYrWzL1CAFpJrpwEpa5aUU3snLpm5dDU
cQ3sIiNpajZjSjGzvotO5CYeQqRal4X0vklbKq9GA1JhpxixDvTNxFKJMySjFtaC0mcJ4xKQ4CTa
gS8QzvDO+pouxqWsE/qkkF20vOkTqk9KLXcJdhXrHG91VD1Llk/JbA6vTLDufQDfs7UkIebHCJ78
ZizNtnZHJeH5CQu2UcR8Z3eaiLowt1u9Vx6mxFApeoOOnpmny6GoovGIXTi2VV8Js60MAiFfQ2dc
9N3XYCIlTxfYaqxU7gzjPWRBEpxb+jmCLibXfXIfKhpwfLBSCDb9d557ZM5haUxNq6hdnlGvsPxE
XC1WaL3WHGE8G22Ft/ajmWRiAYIymvjk3gH4BtdKoMN7TZ1avUBTYVb2bePYjaSWVB0HbIsqr1Qw
AIo3ez8pTYWJzNvCgetD78sV3/GnI8Uh+tCV+I3TvTIOVszvOcObrZSeKl+zHop6Ugqk7HYVl2t8
E0FsQgDIQjUou8INuz9KX8NShlP5w78DGFxHTgcNDKsfmQtPR5iEwv7QCL5XPZ+DI6xvSgBub8fQ
B+P0TLSDj73yhLwH8x0oVP9HZv0x6XKodekdtQ5ZHtVENOYdOaZkZQAjmMWG8soBdktTmXyXMCPZ
g9hmJ0dz3E8KRhld/MlXy+hJ9FVlxYX6PpQcObYB/UgJOhjJ3T769XCHwRaQgNjmovxrfer3P2+h
aWYmxEq3VYjB4QBlsrnRNav1nTYJvWg0ZbbYe/uLUuT0vfxhZ5vd0y0531/4ktb6KRH25gXwDl+W
OyiBZXs8m49KI/+o5w3zJwF/FIHmD+MDPd9ygYD7na/Dpbm4MVVt+8RcBr8JRte1noOhGqOVG2Xl
WuA7/LJIhRg7Uq32wX/qh9QNpgUEMn4+f5V+D64c8fy+9Lbq/3EckD1gTg6qLWsEjgTpXVZBYn6z
TTDZlflxNRwznO272Gme0eMsOFz6cQyv6nHokriUWRQ92Pu0UPO+P+YQkiJRUH/Mx60HSZ8axuu8
ZtXzfL+akuiQ+/fRHQGZzZTGd1/KhtsIPOKEGwGwZWtk4Z39HL3M5mdSy5ugGzKutl8qdk7KY4D3
JMDjcusG0B4IFNUrqbls+S4GFmtDOWDrtXVkaeMOI5HH6+VssSphDSwWYPpZtzfjxDPLtr20og2x
A+trjxghw6T808LjXwEhy8Qhh6MIJhGJd7mZ3p39LY9zp/8u2JgO3knLtMJZzf91BA2TxPVIsQtQ
Rcyc/UIsBjcA+iVNDP02ux/tDARvq2aINRuNPNgPr00psoZYj0pgIqkfY/xou+SuTQR4x6JhHVML
+ugSR4QSDK4udRNzREnYRkcd24iS200EcsI94PolttE0URhOThl2NC9JCJ+iLUBoa3U1ZE+VUV+v
DgX4w/vEx0GIP54W5u358rF05/rgF8PHhrO38jHp3s5hbJuU6jydDkMPK6oFBGesv2DLG9RZsMVU
iRkyrT8+6FsZEWBdpcXjkPIJjQh5mNXycriQRIDTwvBy9W47v+LRHks2O/nUlLHFaXDNVBnjNVTi
Gu3WSuKUYuaMhikdb8E0If6b8TYdIJ8bq77nRsJUlKs0y3uEZXnmZZi4K0UQbforhf51IvF+QsxT
WQOMztfU0RGv+HcOBGZCSLwdmSm4o+gJUcfMioMzIA4g+3EMbdwBUri4KFJwxb372nHOTggP7e5o
9KwtTo7PPxECDeiW8pKlZ4/Vvb5SRPfDEqGRQBWqu+A5sV8WvqZX+4jwlEV9VLKtFUv0MdjDDxo4
xHIlfvgPfMgEX803arURN2Y+kpj96PbtiYPStaUW8DgxsPmGseYIVyDnGT+/XYlQi29uovNaMlxp
ofp5RVtgQtMwy048xiqfwy1U1UMvMfggpdDIyGnW/wJXEsQVb6YoOuxM+kmFFTmaqDzYJ7VfGnd7
lZRmvZVOvBWVZH5SWpCK6NK+sGcYQMYtzUujmf1MmLzIQ4XVDjK2X2zmF1yw5T/V/UvGueICOvFX
XLsS6pVK24tAZFePZTcnak4vnf7oEOFzMjwtNcjQx45bBF+48Wrhp20K0Byi+CO5S7Csb5Tq27OJ
vgHUBg+5OY3sE9Oc6iqd9uhjkJNr5cU/iNCYXJyXAngeXnNmfS7kWR1ZlmrWX8b2j+Mew/E1aHum
SFDDQkbLbdkdN/7CaUlD4qTf9XHSOPqefTZifnJKdmnJeELGrGjIED02ve7ABzuZP1+a3S9CXY5P
mJYuy7ByfbJYu9Z0ttbgCTBDnJx8okgO3UG0aRF0Sf/nf7OGPkC4Y2AsEk4vOKA+Aup/s8mTMOqj
L7DTzCDk31qV0kLzENIYDhBmY+8DRu/q5RmOdsjJCXnNeAxDL4/BBBRfoIvcCz9Gtgp9ghBMWIHb
E7/KoJy/DqWXUm6lS0Byz0W1GDEfOPm1XJuF+C8JtvMQ7H9mLWevR7menRma0WGnyVXKdiQSqOde
BGYhUzWeS79QdYNNTqt41QDhHxg+D9gUS7nkEHD4+0ulpVlu/NNV0UPrXJd48iewb0SOFi1ljOr+
tplATPto8n5CiKokHCAIcwW82XxZXFCgdBqnLzDTl9UXZEdPZ94TxoHDdC7/E+Cf8cIzm21aMWi0
/BBJRUS1Ik8RMWRJrHo59QWQAc5iKvqq1FGGRbgBJM/C8ykDcy9KxYIs6xv7/dTw8ZM2vS9sxKw4
OC8DG0iKEEZGmPtBUX3Jaw/RBTPyd32Aqmu85Z5klB3rRWAsWtW3eI1PWJMUOlzh9A1ge/T6fjYp
Zjp3E9asEQxiZtzVQoui2G65iFtIJkPfZHnG7ncwj0dPgRYvS/vQgFdIQo70Cs2ifWc206wNympe
+HNxoDKzyBJqdEuRglQ4LvKqY1BEyGAXW+pK4R+ERaZL2fFre6TLZfNfJUn/+pamt0ngM9OLNni6
es8CKqQPQmN/pc6O6wKSumodmJzSlf7On6J+uQ3P7K7KbXaZuAFAjj14BVFRaUjB+BIuNNOXkyKd
CkDzf0BULIFqf+X/7j48g+iNfW08uowWKpnL8+jbmnxJiSkycyDhqotiRgp1joE5oNEFePdjf5l9
bZqukDRYwc7zXoyiAqCCBKx35iKmKAW01WupxkGttYZSc/iB9HaMdQV+Fc8cKY9ra3QzFKvvQPFO
aQneBmrBeaS39fOIVRhPvcTd3G40HkKjp7i+g1ShvDW36tEN7F4YJtg8tM3Lf2/XSmxBZA+XdvGE
uM+AXbqSvdKF9xfMMILz5yoY/Ihg5eaJNqXj+8ZIrBsHWAFUkhh+vPeKwkW0IsSjjFgPcoA3j/DU
KipZ0c9EC2q4Q9ycStYBo4sKt3Y/B0eSL8hOOxqSX8gkpW9XoWok7NUXlBI1g+hezmiAiAZov//I
pPsKX9gJpBoOwPndlkjo6OfzGicjOGuVhCnh1PGJk1QLnYLK+d8G1G4cwZArqXU9T8jtUpNDSPJB
wjw87hR4UEKPSRMcO6zgMw0brZiTOKix4BXPjwhup5LNyjyFahhkJI4tdq8SUmmmfjTxBrChP5bU
+jDNDfXmudCOEx1jQMPDmXZfScVtaULY0DUqzBQVHdOGJB+HnUVB88EKY/LPAGVyZIiYg2ySOFKG
wZIICwmVyuLPADChByeaw04lMQvwoagi2EwPV9FklXPJ1tp2SusOZ7EnNNdyWpYLAd8NZIUr85CU
INoooAiz+6ap6A7DxBQ2Qq1wI6hEFzaBBegF0+R1VxAbCgVH+rpl0jwE+QZaeKrcyydLdojnDjfP
Isynkn2tRhgn1zOAGZwYbLVJfI2IQc7vdisWN+ua+jlPs7ITfwVNLcwV0cTBDXUkg0TSiqFNCDMW
yB9Klu/IAv8hlGk3TM6rSSHxMvWAv1e6X5nEkjbD6V9k/h2yHWTZednXT3ON4M0Q5Ca1m1wU4KGW
GDiM4i17c3OMUroP6eCS7i4DNLf2av3URYIf8dtDsNiKYK/6vcpvLJyDmLHeT0WbDVnV6zR7zUBC
jIPu2HtgKVg/GMYJzSo9qxWg0yMzDFVazqXd1xj6kJh4xLS7bugz+JaQXm+G0HDXYjfOlg+bYhXW
HVEKefPiX3RjTca+lPjyWdffZAtr0fU9kb/SpcCtifO97ihr4Soo2GduVPHAIQXMd7qkfpfsX6MF
emXHyOHXvBBC9D/Uo6ChihjFIkhScXnJMkhGAts3vC4eI9L0Mu7BJ1V06nqe1buFSxIuHOUUV4GO
ehFavww+pF4ztPePRTpC284LGX+L0THBjlEkSMv1iviLYbAddVzSAy/gkHAzX7iccDPjnpLNvf3s
cI72C6xIZ4EyutyBd2KVl3kXHerOTvvH9sT8AbR/vw+UNF4u3lzfKsJxFGNHYD9wprOD3cC00l3i
cYblpqIB6XFkq/AbGEPVl/lmPDL8+sUQRRFbzLhf7kV127XSs9VxEF1zvNrC+YnSVok0G7AOO3lb
3ZCytvMdulpb6W6niTYHI+CKSF32S4Ek2nYxTKxzj7+tYTuMbm/30ntDeXK1zB/cVUZqVpgbIalj
ov/GyBi07U5tjDKmipDqxRIEFn71i4LtPquuuRwEe65iX1oSXwU16HWwVjE289rXmu4it3wWrjo0
YhlcMobIIon0zmUbhN2frXuwcC7ovQu1g3ocpf/ueONNwqFLng9GVRek/rHlgkPnoqwF+5C1eV3v
H3ojkAx0pDii79LsvUZ7bqG8E9oQwoZuckzRNjPQ/E5NrjJ3a7mxlJRasCZgYz5Hx/BtZsjcpvvG
2bOHXDmnw65k2M6gTLMtoXx0Uw59B+Qo4Ahgz3M+OypjChwRacmemV2KXucBLTddj1NzE814GC8c
Txof6vKlBkVfsOlCiCyVfomXoyyvfFkH6thWlfQ1tfMY6SyeiEsjd6b6Kx04g+wVvne1BzGoVY3Y
nH5ptliv3m87ollFkZKg0WJkrjAptfx+QXA5btkF0+y46rBjXhkLLImJgyq/mJpY2ZmdsCYqk0dT
SR98LUVfu8lQZDQs1cjxrSG7BVUopMWT2+BRuDyuDdCGnYKQ3m8LiTeAt9/sVSvM6btAPV7ix1ul
AAJdRqCGUx7M7acRQBiCaenLydwIMfciUaJjj8r6zMqErTWnf0LZxTXXWrAIPxPJjv6JiuFp3CNH
6ldONH0DT6PhJNDhdtRPJUp0JBpnDqGvEJWjbNULeCmXIArnCa4o0WMCffhR5kKl0twUEyQ5s07r
DXXLa8xPHdy1HXnDkZNVop3RTfUFYFgHN12lFZFYZhAsnDh/BRpj8lMbo4FqyxFhEXFlG7rj6JSe
ZONLJZfhWIgysiKREb7u+XuFFw9HPCmWn1XB7MyK6Aii/PJuPHtZabNzIu673TJOBYv1b3/FBk+R
y5UMK0JkKhHE8abd6InSD+CtJ4BM9/SROJusq6uLqrfVeV0Om3YFcOOMwmPbbazwL+NlN+hx1fFk
8Y5rQuZLyqlk/OwyH7I05cZFJ8wsS50fIS5Sj3J3NHXNjeCE20kHtIWLyMcAqBQm8n7DOphNjoeW
mC4JZ9YfaVpKxd1UBQyjVPKJ5KY+vOkzl0y8IywnY+MOn9r41af/gzJACjwkGn5TSils3DSp2P9K
qeSvEvfGzwkWqP5pPgnmEfksdZHnq3S++vRLiah9JKUG57aEfSYzKuM6P+b6hcU5WIVIACRWNBqj
JYw8JpRRMiPqwgjC57XBi86PpFBs6rCo1UzwVFeMasHA6qW7+Fk257b9Fwk+IPgq/x66gxufCzFz
8U3AJd5xWh1Yyq0nB7KE4jDcPaDqgs0hDnj8c3L7c+pvdR6EHN8l6WcPIZnp2nOsdA5aH2uIYCoR
m8kk09kpvmPbLvg4BOzFCDDoK3alRdarmDuQMD41AkJ5Nq5lwgJpYxWE8xaWbnuWdpgXn1iJIgug
0Mj75TtWLizMs6NgosUrKFLVdSvVF91jEHa0HcmoyhkmUfLHs5dKkkemAR8d1jrTbHYOcNEn/phH
594yBxdOiw7B3G8qj+8Vd2CqbXxhII33SjtbW6tGviQffeYOj66+UH/5dxXo9r/uVrGrAq0niFju
i+s14VIlxBOAszlem15lk4kuU1NMralWOm3AVMaBBRkkE22V9tUpe9Z7ENtOcwVO6ADYPGHhX0c/
qJgIQUpA/avEz827sJd+dsKeLF/5IS38Kjks56uYi8KbxzNs4OOvmF3717oN1P7iy1tcXHZ1n6JJ
zYppJmOBSu2XOgLTsqWpvaaAxGVGySRUowy+7bFdDtfJE7ZDCEnFKdCx+5gQJ0lwgSIhFzlYyWHL
2jWnbfvTZpnHJWdO+lTlmjpIJkmt1aNHlcIoKuRYjbGhfu+YFnD8NrVeWzvW2LXj8Zmj5AH9pgrB
CaOobiir5E7KPD8m9XWqE71HHguUG9zfR7ZeTZU/F37Hhyhu2Z+CRGB8n+7gco6zyZoCCbk/blQh
yVX0OyYHw+bYxJtjr24UWSsN1QuY4caSFfgB2yg4YOpLIAHHiix8ndBzk2oKN67zvcWdMrh6myNp
Hns7oEVzl6CwhBdww2O+I9EL+JfRNLjf0ss70qm3FKe14ZLnDVNEu5L7pkX83E5wbMQLoDHp7nfq
e72le4/jy4bRW5+bMDmkCYYy8HXGFGEapBZKS1Lvhs+phxMItYdC2Z8GYL6vk9P3OY2lgZITj88o
fkxwbok4Ni1wzwAWS7P3k8fxORTdgW8pJCsKnYQyzPw7dLGHC20OdLdvh/aOxoakeh5KmsLA1LNs
XZwrMH448XY4lXX088AmiHFtcf1Ju/dJeHMlTUuG29pWc7exkfYLME347Xgt3GWNmsQGYO4WF66E
SJmSv1VD0cylpdJUdcfS72oKa0M6BhalOdWZQShZK+WuMkG+6+oh///ZJM16goavbbazqu3oPVcS
M47+IaoQusycyGxTZDqiM3oaZyJiRGy++1CvRIDAx97LiugrMK1EMpqJKfnbzMkEyT4kdVPCf1JQ
nfTvpgrWrC5qJNWXxAmRZFrBfBNd1MX5EtOkUnNrNpMHT0TqvCJ5liHKdcZUh/LSe5x5t0T7Vnr5
T4iGOW6W8sleburc6H2UMvwe9vuPUzyu+WDwiRYgrKmiwOaIyQqMzzYudT8s5zrnucsHmXKEEa6u
c7jwrgKD+YtFt7vHICFLuQUA+1Fl2Cog3KtFjVq+6Fi21DwUW2DXwioc5TpAj9xZG8CuCD0gmNER
+2GI4gSQli8ThQPNXBN8e7mDutgRfAdF6KPdlMjdE323TVP8dJm3Tzr3zSNaVuwD+QS9rpKGmbRG
QAI36nLBtfFLYa3IjBHzztEjj7jr0K2gKskJPCBarJy3WKDQGVNPrPlHLyoJnqnIxmWjCgGPENlp
xd6Zfm+WzK6pGKmyNZtxO0C1V9wLG2WJFemGJpX/srbSh7wwvdtm+kk8J6crC9MSXPk1or7iDxhH
nnTlSdnsb0btFlgPULQLVyihGkwmO9yljLfJBFU073LSWwl1urjqlVM+bbpkF56Yi+CaKwL+ZPri
blHD+z3mwbkaCEIIUENXn9RHkhfWuQVByeZ45rvClzpbgDQOpxqx4lOQzKi146gbFSFaEVeZQSWX
0WnAG4AX/XsoFZrOHEM9bUaaXJSmqqxLAelsZStOyXqpiwIDgSi40J+V3mgMwqlfpKrBxFOjdTIv
pCJ14sHxrJac6NYDBwlwqOhQL6AJFQk+ORefR68ecloadr4RlICo07F9TdHvVsPpR6bU8WUUVGcJ
jJCh52p/rPtTRw4tigqDwb6RO7wwt+4bzw7w6aLTswZ8Lbntaa91g5oeMEyS88lZ57/kXozel5he
K0ZxbymLDOozFu3DszuNeiiFS7/g/8dSYWMlZ+hMDM1bmkw4Hx/n61S4UeRRB7ZR7ehdvsjTA7Ji
gdWpnfgz6DrH3VOJzc6FO8kOwwEXeKhcMOTyTK4DkAnGLTqL4fxuWvfRq2jtAe8BeacsCuNbgKm1
MWN9GK7SV3wibYsDWgbkYf8Ky3XBbuiihCa/qddYi/oLJP4TP8WpMrQlJnT1b8hxf9XSDlpneyX2
fsm181qU6Z4TKVJclWWbNhOeQnXfg+dYH8sJDqpzOeLRkbhf+JBo0zb13ZggSySavNAwlilRZTYk
fWlrQZqAhhDwBJxR2HjO75qwSTCs0z8HgYhkSQ5TvXhBkV2qvUfTW00X8ohaIvDhzPcEdd7IJxhn
xY3VCKn147ote7Pwjdv7OHJLYp+mUHhm/NsQ1vpdQEroMT5VPSfVkzvRsCsy3C+N3YRmLb99X3lE
F5BeJWZ1LEs/R94bcm2iQlR5t2Zwkkk/E7NPPfrYENirpS9DohQWw5LriaHYwCYvTi9dtGIUp17P
UIl7qFbCUNfvwwJSyruHwJe26wk7ZuV8iP5+x0pePZ+eYtMpY+mAEqzzBoWm7n93ziQ7BcurWIg6
2th3glHNXobzdDvm7FIY2f+DH9/SDrxZyr2AIN9Z0ObeVQproy3bQF1LVNEJ2doTl9p+Wz3sUwIB
aITkfNh1aAe+TCDE5A1YTb4Z4ZS+9BmqZ2F5pMRH3qqBMa936dH37hnjz4a7gTW4gJa/e8pp4JKd
2XtwgIXqulm5JC4R8DHriL804F6hrhnvN2SjeX/1FRaSAAOPmSv1xdHJRI3Me+NfHhaUOUEcH4oV
pBzfyLdVjflxHU6Eau6ksXvkMCQ2l65Cvi0uLQJT5eTQAsaVCulBD9Xd/nzYnjEx/YSZX371hFOu
5nHSwjd45/vqj3kbHCxcDDP+X52/bpK4Hs9GDERcVamrKBZEL+Iv+RVUG97RDcbyLULz/kpGQ5es
pdvjbWq0KjjcsEqTQ+nOsXpPZhen1AwXmlJnWtYct77RO2lxhDzWoUaAs7y1EJNT0FheAhU+/kvb
9t/TLfjM5yqnKN4qgmXMPKXacX+ialRxJsLap7UYoCDj1v0aJgHs6HTjdDUyPMwYJIeRuPbk4S57
NWBNZ3LPn5J9GQ8hioYwtv0Y22fmKaSQdLOac7YWuuJx28eqTU4hG3WlYcwVzMGIATXsHYluCitr
NV4GBQkGomR+eJ0tikZBwWY03BsdMQazyQQNjPWKMRLif0dHWFaBAWWsm2PWHeppUC5fmhDaAwrT
yUmxPWVo6JBk+pQlNMWKJU2aHqfygsHGZX0ICS8k6rlYIZP5nl7VoydLZ2J62iT3jlEMnGN5PjX9
pC6DwAMo7FweKydZBdCedGuNJhF9i1xY8L/GAFYHeBMQ6LrSfg8ShYP5dzUSOXT5v2n5G2JH+afl
Mc6ztX+S1kfbxOp5ILndjAnIpdfeNm1h1e0u3BmqBmVy20PPEa5W5xRWLrRIVBtuBueD5sYAwVbq
F497bAkoP9fXC9BASzdniKkKjy8vZzjhChgfyz5aY7akyIKb24q31RkJf9n98H7+j1taoGrU0nRq
5yrYtUaCFPHZMfZJQYgvAF+yRW9CqBDk2TKa4O80OWQcIEZDAUJdr7xc/snv95+RuuCf/pUNSZz6
OwrrNLmtPU4epckgwt1tfMySoXLsX1pBJ1vkHiaewqlhGqwdr85S2ZAAG0JfzwabycOOMkGlAj73
WLiBhs6kRJS0aP9/q+lCMsPx8ZFO0Ceoe+a+RWv++5e4dV4hkWudGmTbYpEmboIFJKPbyq8OY2R3
8PvSoF0kaOxWcALpX6j8iPXopxD3Gtd+14QCW9NrHzKQ3PsIb4vH33L4hMyvGCC59Y4N4IUJilHd
mtqzOIPTLEJeqtkLZbhWaOszYCra4U5/H4beOh2g0p6+ZaqC0Y2V3godWq3AL3RAAQCSvFrQ71Tp
I0TwMDAGk/cRSP26+V4hSIAFV0molrtFqRaaZET18Y9KBqW9tA++hyrCfmI5U22FYZw9yWbtRz7A
VQtuBzdy5s5F5Z5iQAj7RL1dVZP3s/8D383dleqlYSUy3JyImC+NE7w+hfX8Nz2AR58h0gHCEnfO
g6WcnWkVFiRQZPd9Gf1OfveviQr6NbaSTtXzRFVF8H+B0oJf3QRnxJKAzuLBOmotnceKndgz2nEI
5MHT09eLv9697PrHIUnxzA5XLq/IpXd7MIcSFoR44AePfYgsM+0FNk8DAPoc0diLdwl44FpUq6ZJ
fzlOjCJMiKYFhHhJdH3m1N1THQeQtzbHga3PnmG+qiqSaga+xtwcOMnW4nkjL8tIIzNPgBqLAr3V
vKWy04YEXGFRiiQe+BFHHxjmcZdUlbOoXTtgnEH7QLD9CgxyrsBFiEcqa/STjjGLEX2n4iTtaBql
/xHhdHsk/JBz8Cc+DkxvQrl9ezyDQrjkR+R1lqHFdkhb1y56mazcxpFBjZrzz0oGogW1HsaWSt+5
rsVnH3Nsy3VF/Dhiwg1Sc+vmnEjcU6Y2+dnZ1vrw0DfTjkTRkK3na2XgeYcGZcvk7e9VyFjzlXJq
d/F9QmX8S7Rq3PXSXWFiNbCc/W+y02I54ohkPyCswOIq4zH46PsicP/BsYmSztWOaYA48WSTRNDI
NkCKPjs8sZreYkAVLtm4IVYoo70hfcCOUCZ5M2EcCddV+63AVaRGGk0oEeH83won0Kk/92dXXBBn
LZfcfvHhylNOIgcYzfQIIhXVJtgbxtYk48jpPN4KKXyVNokOW4bnufsmjsuP9Q7Q3EYtal8xie2R
r4gjH3cuIIsMJBPtXyX2WrjaS3+L7tLp0l+RglHBsUi+Itl5kOJUdZw+AW40a8fmV4D9+hkijCqE
vNUxp2VH2VjkxIjOhCegjrpAcpVHLW9SSx830qfXcNYOs+miBoInalvOpNr6tDfoWeJhgVu4VEQX
1NFXitrrAh3B1sUJ4rg9wvSpoWBEmLlsE60MRKfaI/DHSTJ5IK6+b0GD43YwJw4EHWA9DGP8BVa6
3DVJ3nLuxKVU21nI73bUp9zNoG5JcbiFR51Ow/TQmfo+T7kqGGh6MLQlpG2+n6wV98obDQNfpPrx
DKc8EO5g+4LQTHINjKMYIJh3F1xPvmDcvDTeBjiwfyslEvCpXRKgwSuFvuSzcW06fONgHpIsjwWA
/v0Y1VEbaj+tDHPxwqQRCp9Bk4qWyFXiEoCyrjBC8jtkcpugUVI8ZmzNwQZowsWQjp9L7umV+F2H
TOGL92kqcWabgk/27T3No53p9oPJMCULK0oKWrghq6ygasm/NwUMoENMqYa12/qk4HP2ithTfelH
+UORODMDsC4/0/ixfAfc4p8vaif/OwMUiKzrrUTbno4l+FPAVerxu2Mt50RRFsk4T808bq7fKInf
X0VXm4toao5AgVAtdF3SC8AjstVYpVdfYnbNk0TnDOd17sQ8ThRogHgdEX+uSJ5LMlifJjM4Hj7d
IaBGV93EVtbReOrI63z7kkbqGOYRtpIMKWVe4+WwLzI6E0brDyCuwsPsYbB9NykcszcLJ/Dr87k0
73dLefxFYPkOX2jVM1wwCgOI6TIH6IMHmF0rp+xZ/M/f7XCUSEoXbeNsuhi/gv5C46mSEU+Uk+hW
L4G15y2gflsWrlsJtQ7KrDqKEqcQtolgYsjF6n3jQy4ppmZkojPtYMSowkhWcZAcTV8SDEbhgsFT
DlVjeyY6zsCxny9VlQ9M643kNo+MjjEkLyUHoKZKAkj8/sGxnQIn9S0sSAq0x5CkuDG6zyQlzG+4
mEuS8I7YyYkQRKnGQq0h1uQJJqCnl5QDNG1RPwT+dSCxTVwUyPECYta5iKJVy0GCA3SfhS0wRkIE
mOxPccOqkUaa1u9Jt6r3DqIPdUxoM9QNOhUh7AMaeaD0DSA/Wx80/faWoFT+vZ7LtKIqsgMz7Cjf
S4G45eddA8vqKsUirH67IXT9MPShttMaQzd7ZNw8UmlyV7jYZ6B/gJd74yfZszt067Nto0pRc8Qp
Z/oAttEFS/yTvus8uHw1lBlsGkK1Aw4s3Ma2CU42MHYarCgBt00XC2WQ2BzTuJK0eHQUxFQRuPrR
4EaUNAFTWubHl12kMxu1A97OwgCKjQFdZWMMzWOd4f1WUGHOQKDCFgr9q12J/65ID6BSUI7QK2hx
zKBMxJMG6p7h5kyc4i2C+9euhWLKwJSfJCwH+ws1RBVPyXiLBLELvXA07kXOvch0xn6ACAKICzDF
rzl3imhb95WsPdPW8+qP2aKVazEfGA+W/YDexAO58ApR0+/qLvlNYEj3OfMAgqU7bHmtXtP0jKs3
+baBbMKWeWgNtGKFcZQ5KdNZyqXbW4hRm9FDVZe2XwM2IiQlPluhkx6YTQyjUlxvltaWFFtsLSUw
hhuSEBeh/j2zb9eKTrskNCBMoLBT7MPLj+TpJEy32tG9KrPiWgcXfMXPmDp2x7Bje9A7cZ8ke6xb
a7G2LIzw49gT5NZBU6K6Bw0JLwP/Es6SgcGPCl/NPVHIfhfl+NlmDwR0g9q3l8WN99oU12cinzfb
FdvW2O89XyVVfHmM9Uxa0ZLrSd/jk9v4vwk9zG3gZLKOCYRx9e/0TYIm+9x8PEMaZ6JQT0zIJThj
zjWZdzyj9gB+qvv94Hwv9CUp00DmAWzfKdqGopffHuigAP1UdCpR/0Ik4NxAWOh/fiWTyZHcTTUG
6eTNd0+k2CIQMrej+yZz1a9NpFPrWBki4QqiIJXh2aBpspE8zhiuU6Ebd7R3kEQ/foY7hpPNcrwu
/6RN4Xci5Rq6EM/4b4Yd8G3eSMZKIFPNN04IF76VCh2kV05/E6GgRI/1+XsKz0yULiFqZgOUmjKN
52Po4GtncWWQ61orxGuy19dalH3InGtyX8tLy8a8r0TEvXAkpNtiohON2Hkj6SYKAfShXwF82ljY
mi0458fAsVxRhBRXTl1klTqms1l8e/HkzKVUR/ftYWZ/r4OqdsiOOqNC55/nV2chsDhyGWVWNbuA
1318UMz6AcWgYZc5oMxKLf7lY0YVxwpteAtijFghdJHWoN48Adeq711ioqc9RHdwJsItNMp3zQcJ
v8L7oljl/L5cvsnU8lw/L6X7EW2kaoSFE/GrbNbHQXo/ZzSvmiBcQmSAcGrGx97oJuCdIRGdEEKs
O5HAhC9PXGq3WKf2ByjiyiXzjDYCW/zg71noIG9yPfhUtcceLmLSllgPJ3V1VyiC7P5qRs/CvZkR
0WXjtTE5ngfxgsT+iOH1cHFUzhVVjNJHlM6piMm8t4BMHKZbZu45V9k/OIF2SpU7ugF2kg/GLOG+
KbTgTPXUMREpnuBb216r3pgc5twU1Bo6f7xeNEWfSWCHaN4qaQEGc7vCo9lpwkoCfd2dGyTFff3Y
9ULsRrb6LlWXCPAO4C8NQXqQoq4mFHENilmDKhYOIyxlrmgQwIrRSQRfzQ3IEINuNWMSNuAdlivI
URUCLPWmRQe6UGUVaaAJ9PWMXqSxxxfiucCN6EQaWHJ99K3soco7tXIP5b9u+iOzCMLPxFg1nAPI
nbRMO4as055c3nug7Oxpt5ZphU6Heh7R/nIyxgZgEE0t6lQyYYLAhq587wHeQW8xvfxg70XjOV4D
YXNIAXKyuwTUTGbjW351NcE4T48Qj/YoCzu/9s2F3QbooM6kKj4/Rxavxl31Z0CFst6ELvd5Dmff
8myq8RQ4SH8Zv5ljuvS1ege4vig6hsI4QMheGWvFEnPDY7iOKSU33Eb4gnnagLKXUF83A05z4sjw
2pOuqxlmn4Cgm294csTeqRvL+do5reJaj/vI7Aki84bDAxR5KEDN3YESLO6lrEybCeKBR+MZJmYk
ipm5ZQfyaAFjVecKoFZ9DdWmS4FVW9jO1NRWxSya9+SOngu0GLeOEkOHzfRl1DfLb8/9Jip1Mz/H
n00QyCbra76No3NjmiSQRuOUbEvBXsPLnQDbxu25BzoUPFw/WsRb9OZw/IQfGnb7+2TutHAZTLjO
vBEak2A3yd7CN4nVkdd/KoTTxH4m5Kvf3CKffh7/MHu5cO2QsdIxQ5frgLc11Eq9yii38gSvDUUc
bmWvqGSDC2yGRGaP6PmpM6Hvkc+B0nMSDCGOzOgG4JXtv1+nuU7AQQhgJNj99awwyx4LYqzHeR6X
K7kOGBufv4bGLo/Tu9aPsbYmR38dJZ7HKZW1Lw6y3wX/8UK/qscFfC+NN1ZMbjtG4tHK7NhO3FH7
yP1N/9YS+DansLh4SKCsRpiFLBCwdLzygjCB9vs2jv2cuBiq5Q+ZQwnitQa+RAR0FOiuF/9wwj/7
QC4Mxyw4Xr7wZrZQDrhhPdhGyDTGOiyNz3EaTlzhkMFVuH8ARh2eblPYRfC42GpgRqDpNKb0r6kQ
EC8Iq20QR8cQsqkemrEIo//6oZRjqOfJ9QDGEKuNNznqdzI+v9LLcohOZlVV2El6WLbGNlqkTTS3
xJrbTq0iOU7YTlPipz6zdLsbYeRdw72vXdm4UnofR+o7pCe6aFgMk/yD7aas0OT8x1Dwi85GlYZ6
UfDpbaI9APbi2sveM8ztr1m3H9Ua+hqKPXb4+yuD0I1n1y39HHTXzIdi06kzBn9FC9M/JCCmVtQ3
tLlvh0VCJtCaih6RvbtPLhXgZu5JLxSDoriKsZmUwY2hGJf43pjqwfegD2LIpcSTqFNZfw8Hsd2g
LxGUqZp8xyLygl1c0xekggpOcMu8/xrnklFTbg8vQWF6hiF/GnOpaQ/ewmJaZJ0dCjNubzmptW4S
4wbS9ptjU9cvb8wqTVdgE4/CzmbbDYXC4jcsPSOvwTeloHGWCO/KzfEOm7X3658EzoiasvBq9cnl
dMLGME3T86gWgqH7ZfkfeJEfAZbxuHhLSmP+xypSVUXnuWMSmIB8wTz8qHDH/PnduKT8j/5ItknD
28Gi1uNfYRjZyN4OMiaRVzqj1dargNM386oiQRZHDtz0qp7taaiGvypKYlkjAVrN9HZ2v2nCAM6K
OuQykuxbulcRGnL69P2F2XGdTyj76TqHgoaL8orMMgOdJsacN4o2EXpTv4mXkkbH6XPDM9Qfk4sO
rZAL9K+6UB+ayw/WepAEW6y4RL2ERRSRCLmHS/Ip5psAa8mOodOmQVik8Dau3X1QWt+oBAD4+Hjq
sEldpUObIyOnV70NeEAguVYlo5BI/yYAD7M9SGWqGIqqvQDUZKaFcLXQqkK9Qj6AHidf9JGDbcWv
VBol2C6lne3uhlDhqpc2+fSMAhesb9PDLTD9n6HwAjlj9fXJsX27n/xnm6jW6pfg0rkaBMoKguif
09FPrXwpyr9sO3H1YIngildX5Wi8spQJSpnJJcJ06sCYfRueKFfizd6/nXz5wJJJV7bRF9v2Y855
mGPRz0lcVaYAUYlzOFsOlCMxvIoiZ+U5W3alxxkUSYhuJybEUHryK7Le9wawXcuIOwQtEPh638TQ
dPdD+cIsP3XtJHy8ZSprxOyD6OiflAlFdejgJ/WZyevjdlLj+3bm8g6ZRpvR8wnPbgQJ/WTAcYyj
CHpHhKnEADJ4n18OnDOWmBOcy0184pPlln5cJweBv9lK68ginUHMYZ4HUuyp6NbKe3dE+FDkV7d7
33NoK75PaWKgLVBw3IhGAYrNHRH2uVUWK+tyKmYqZbzwzlq5CLyGfA3V1FB8wnLko0kWI8nEog+c
cfWiPOsX3vCvZKcJkUUw/XMkCMRJoMi7QbbYykwBJGDDiFoSYa264i2vl0B0JPuKz4xhWPBxsHK3
SyIuVKsu+Cbp5tOUn6ThvZ0KJ1ZDh7Wk2rdKrb1axcIzeiEU9eGqccOG9Pt6fhejRFVEIqdtkqNw
+lSPcB9AKUDE1cMgOvsBcmyOeVZToDdHz0ETarbQclxf7y4NoK8YzXCFZhpyCmQRPXCMfak7TWRr
2Vdu1WTt6+YP+6x7umr0lQ35rhK+yNwCltfYL7+oGTdhLpIYSz8zg8AKcKaiXK+BHHrdpuaAmSGV
TqGXwjszxv29c8zaWzdQzOSqGE++9LWVCHysRQSmGdyi5fcxbMnf5sQOeP8sr3PJO7jI7YNqUBF+
Kj+U2j0q/sEeztOj0eLGGe7EGshJNPlpKB+6bNe6I7n1EMNuBKgkkhCRiufJMSSiXzq0L+JeHTLj
5v0aTN2HuP2Qqgz/jlYlT2KT89vm6cdm38QpV82VfIsX2F5IE6skJO0RUfVD0/eGn5GjcOFDM9Kx
c5QCjdHLm8Nf0OqGrLH6lOBkV8+hR68yEhG5img7IIq0LDfiIZYO8fFwgC77AhLF/zm3VvKOBXu+
ai5vbZyc2rVDY9mRPbvEhEs81FRAMaF5bYRpHMTBJvgQST0xvu+Z0qVnjn1S0vrkUx1C0+dzk5a0
Reru44WDqGkjTf49/TUC9XUpuSoELYK25oCNDzpp16sjSzAlfQSuXh9bC0d7d52eotQc7q1IANHO
4hfYg9+GA1XoqHTItZ3rq+88VNz+cAEIIsBeNm36sJRStpsp5H54tHCsEGglPAZPiGqx224UwPcO
FZVzBOFaQmMq3zjyFcJ29dwnDDoDXa/I7WNhZjZFby0DaFD5h8GZbZdKRqnxKPvN/sQp7FhlcqQ6
cfU6JRLXcVpl3qf7O4GPaPwOGmDNY850dTS4lC3Y8177wf7ymGxkXzzbTssC9bwYYXTgvQQlPAp6
Zqk1zNaOgSRiJjbZ0e31GgRfYW8aoGORJBkMZEd1mDypK3YFlVc0bYDDMfsOk8TIcmDD3YzEckyk
qpYsa4phOmJoabwyvrWj/XHIIqrbwlePJbIzm+j/xdABkoEpehXI6dowSxIOPgkAsL0iV/3/BRmX
wxpL0AfntjX2qGgGYgMNBC5awg/dW31mj1Xp7N7dYLTgaonqGvhPnupq0Nrn3MeOuxzrjJASPdzP
AoeIlKURnkUhRI6TpHcu20BrSwVwnZg4ecJnuLkATh1tb1NX5DC4jH/CyQyeBZkcoAIOpJtEKQck
fJ0UbsGSqKZ7YKHbFVhHRyzq0g002J2TVOiXYEA1f+sipM6Bvs5HqCa+ymgDr8fQEGXP329G7sZn
qnh2UEBnrakjja0WECWZp2G60zZ/YCsj9Zi06M+K4L7/yamhDkuyT/1F/QuF00x+qF4c/EyDZvvX
BuT7a2yEtq/Onf9/4e9NSQc8YKv2cSKd3Q57WBRbodEiRw5kZC7ycCzlEUNbafZbYuAEaoNZ45gL
7QSr3WjmckMNI9YsHQtKbB6AMEgOYpsnIN9dNb8MNb+oz0JaggqRY/ah1jh0B/HaTrye/9jAJmnG
EVtEV3AEi7qM2VKhj+UqfFPiW+1pZlUyBkSJWBmx7G6cffPMpllc+aNV0aIJ/b4TBrIFpqmOTWsf
SHxNTCfP1w373MEHH1B7hfVU8ZJ1F4TjVZNoROKeZHc7FmzZ7cmVn+F0Fqji2r3onIKUM+qXCFo7
PQ6f+7YgD3KiylV+0xgP62eRzFxnFC8j8dyU32xYNd630plBiogAir5ZXcSjnTzMkHhpbkpG/oPA
sjVMfmXk0dveCIA/iVTpe/9K7OrlL6fCsEMZ1oQufEyWiVB9ErR3P5pw77EdS3XBgCx8tpvBWR+O
+cvH4ZXmWB7H+DIfB2maGC0DupgdfAC8Nn1GeCXJu17Vpei8nzjcd/Q0vnHr44a8nNdJKxA0PbYB
GJIIcmbxARoObEE4G9c1ceKCZalzO7fozqTXLma88JBNW8OHK0vR/SVX4WABOvaa4lfqbSRrFEFH
ss5rGcUMt6mkrnUVzwgEAnu5iqaWXVOv8pwJ+98qHd+ohWg8Q3SI13o+IHiooEPXw2NN1KskkWtG
7cc28IWfIGZ7fbSG/yLv7vYlB2xdsWACFQZMEsho2oG0QQkneKXYTdnScbjp7zDbfT7KjRhIPZo4
dAME9p1jSkm49BXnOiz83ZfALjdc35NPzwEVAmrJw7u+OXSye/1dHagqKntHl2ppBqicmZgo1OOc
tlXlQaqj5BZazNdVIrCTIj2aNKOkt+mEAjSDHE9LUONPaS7H48r3/v52vhZOQKwcOcSBI3YVYsbg
0MBpKJ8Vsgfnvz1NG6biXzVvsD6vYl/H43WTynv5M7sajJq1EFS0Ixqa/Q+x/zjchOqFWQSoiPSi
FQ2EWUyesU4M6UXjMyTbm0GOb+wopmk9Ub9P/TbWdyQbKGuhj+XZj+tSQb55F4zjBaUKlRyidVVL
uGtW0SJ6/CdRzTSK40z1T6+efLL4lg7LBS40QhoTwWqbbHuQ1tFFymE7OBrVYN8OAwlVHJ/873uo
6P/fad8hwR6Asc9SQMOxD818aUtLSadjzDJ13aQHJnjsn8ZOiEwkR8+Q0GpPEVmygDo3UtuoJIpA
G8stuws09k2aqnAZ+gdckV+OCLKoPzonbhF8dfqFNqxKRow/LrIMzhTcy3QxvVvlOGT0GBeS4R53
rmlnK6FWXoCxr0txYLSdsUw5I0QcHF6icIW9pWlrzKu9g2Y7EZO4TL7SKRFNd/Tg7ERNxBhS4rYg
0b6X+4memgE7hA8Xs+CViSZoH0/PUCgFvN14S7o7d1mOk1PEzrTWvFTjL4kRD7ChStdG3IPS6yFN
lE1UFi0JxmQ7yjayrEnZTCPmMNIemKTVgYd/i11q0zHkegeiCpgadcei7cFIM4raRY3oRMX0sR58
w7sirSUWVRmKacSw8JsMzyqaJ00ykbUczjWdhhUsKszSfG+gCFR0DoH2574lE+YWiIzMa+VgCJxu
UfxV9rhJnNAlOu6jpD7fgWsjgqPQT7X6DWZqQ6Bcq9do9HqenM13AUH4sulzGqtle/kJJYHgWsz1
CtQ68pooVA5rGkr/zjY/kX5MYfvzZMvXLJtoQXOJmKtRX/UJjGGyK4T3yWk4AqbxKDIk4M4lBTCi
oShKz3SjSnytdBET0hm+JftooOTKu09/z+wO+vxR1PvTDlxwIFTDlMr/JBOVE1tpGsA08/jOCadp
xdpyYwzs7ScsHYPWUxr34yNuGX7YpAGi1OCQUvBCxr0xK+4kaM2k79jp7DR9r9c31RAmkd19oYDS
K5XSO91ypa6TYya1Ld8/V0Fue4eu/6s1Rh41H6WT/BoqCsHp+6TwrGiOTDAXs6UTEBlskXiz6087
FBCbsoyOjhF5/Mm6mPpUhT8wJcrAasHysreppDQVk+EQuCXd8ubNf3L389b01NS0FpHw4cwPVzaO
HesEhp075M5tqRla58YrLZl/7AHn7XtOqXZ1RtM09K1wZB2SsPWdjkWSlzrfi2KyCYp8u8eSX+yL
V3kUB4pRyjr9OwV/mKoedspQaeDcnYaMOr6rt50XYKMgp46Le7byO9Ru3Sot9Lg9IEiG+bSH5BrJ
iyNKTFQEC4jj18ztI0oBuMbZJTWZJbrVGY/FXoOYFcq9Bt/sHBKoP+Oe2e+p6fHKmom1jnqTvr3Y
lEJU2vaq+rIY4wa3BQh7eKmUW42+EoHOTsozzMwEcEigIk/Hg4EVALwwrZXatvyaRnT0O3fmRmII
E46W+3UwQEW8S7Cr8t6VfXTvpPpUV40Psrtnk+itj41gC4o+zmeiwKoTj+thy71VUUgwukIjhNXq
YoYgszMg1l0ePZgkxXhhg/RctEh4aLumd2giwHeOtQxJR7SJz1IK+bmgW+tPzd+vvAJhmU1LCM8Y
igJVjW5S5KAYgeP3xBzRSRKDt3rTXIsU41EXHQjmYO8YsJfur61lDHmkCjF35gABvvSCgBKoTgm3
kO4IMG6x4yCxcklkrgFGfTNSrhfezvt3MCjxrlo8M/upV/EmDHkQgGNgxrq8BEKbhbjX35WWm5K9
wWhEP/E1fXJMOH1+iA2htMcgK5X0wnbeOp8l12dGJWu2nnlVqMzaaiwHkDD6IVwVOxP34/NDOEKj
KbedVKJwNJjpx65zD6ovTivs6FQqri5/sK70c1OVQCmNIm2N6sKVQF2052ypkJ2Y8oV4PO0lnW+/
A0GpU70dr+16VjvkqbXKuniug17Ie3Ihyc7iUoPw6LMkzAHwkG09gTAQA94+j30mZGvkNX3KWLuO
WyWssk9EPFAWM00XyQmMI93zxay2Aqtz3XwEgcMO+n+BhA3rAVt77BmwW+mT/gUkMjJv2JseKiwQ
0uWaw7W9b79vkeZX3Rr1Il05fJadTU5Z9oo/YaAcRIJusiqwZqKLKn7blcmfq9E9wzhzbVpdK92d
ieHe5k6JJEayyNvUEpFv4qLBhBNJ0EaApert5/P14rXqJkKnqryuaLh2VArS1kdsC9BnoKt6o50i
YlQzUZDkrwzYFgO0IAUP2kUnrcnUx9UsHnjkY3d8BoLTfcgjA/TsxDftSZt+z/5wdwcxDG8qNFD4
JtfV/afv1ZciReAZDNndjn49D7r9nzsvUHJ5r2NCqAUPHpNR+QVk0Y101sTSjEg+NokatUsZBsDV
L2jFuH2xkP5wBX89t25Y5kOCVpxAYm6oVHOkzAFlxW/zyZWg0N0JxkOZIQxHBSP3X5fALHObyj1Q
CBYqQRPN0UDwDWQLoylSvYJpiz/4spspapBBSgA2hcZBRRFIPHqVD9R/9G0FuuCp0rrY1znclrHi
4qd/bjuvdBWMPJlQ7CpPYKW/yNIXCqFqEXL3pHAEsGomv1diksbKNoyBfDiyLi6ATl+m7+35a5FU
rK60V06cVyn8qnitvxzbNZ7lyNpRAAJ5t7qa1Guyxcifc4Iwd8BTlhGrdN9n0r3pNcAKUv1vjY7o
UQAULHYI8zkmSU+dBgDEOWOURrSVP/fl4GU8xfkHjB1b2pgG07iXxkWV7fcKhCilFNgd6kiTGgtN
RWqf5LbTa/j7FJu2iG4TtzDwnjY9Y4mhALbKCejrlB9YQXrWuzo58HAIk8uIflplttuFb1zVM4dG
jS4ScY3XeTJJnF93TaQDvDJWT/buI/JrBKG98fgFYQKChVVXPsHC58A4Jp02KPE4F6bZVV3uo1LE
pcLTWuXxaewsEu6/lQVrIbfCJZKMdWnfV7ZtO/ddkhlUQxBzZdiqK8Ms/yloZLOGs1Kpa2irsDlA
9VDJjs/jLTybkAOfce6wNLM5BM2JHdYcffRWtN5cqRbX9Yz6pEb3ztnTpUCthC8vBieVL6M5+81q
+Yzgm7g53/EitdRNO1o/LeSlB6nubh9Xl4qm/O9jn5o+vvzque2TAlyodZ1PEFUMjutbj+qvuyWZ
mUuMMlg3dd4kBiiuXWsr/8tacFQ6BciTQEkcWLsT7wulXPVPzUxumZGYETMr53gBZ+N5eIGM3/Y1
IOFg3KvlHw0JUJOVDZkqWJb5HJlnJ41DEC86UjTvpjHufla2qdbF07a7nv5ONDq49qf3VWyQ7TD1
4rTe70rvDrw1h/Mjt7C8oytto/P2GCNouueq2vgq7E+XMb5joUSFDqa7o/YMwgJlNg6O8U6O7aSm
QGPExBlq7hfypVxYiEI7+iEFQy0I3QcSKqGjYVrLwYDCDXPTQ4A/JN+Pv6dwdk9g2SHK6nHm5LwV
wcQmW8ObnT8hkxgw0ZG3EJsWLYGoHJ3IKuM9iE4c4H84+6modiT6TShefBHSbjs6SLXau3Mt+yED
YnF5GJv1NTxZ9AePRo/9JEfszUWM2lrrd35KsBfuH1kqISW0nKadsS0yf+Gi4w1e8VEPn9dxnaiW
Xt/t0hstzTKXrq34x1D1sOWKTIr3FEo9VGbQ8Ah1UEUoLikF8KrW6AYCoFgy5v6M2zhpBsyRYqon
Xpn0R7cphFOV1V3yS/mR5EOOhP40I+EABO09Lx1KLrqcMrVnEbVi8whsbLaghvs2Tweik0HtOCGV
dNgzGDJ1BMdoR7s5tdjqYV+jJpDrx/3yjZhXEMqyBa7QGbIs6/giKDF3k/MTCTgJOey925mt6YtV
0UYJapN6Z0jsARIuRh3n8klBHHMlXU+sSVB7ljHdznV9psMuww3L/waC+lMcQkhIWyV+Bq5/Sea5
uD3hTBlu/SS0h6C6pzWiUXgN1FN8r3FzWl1IhBVYIbgnMrpyvarXySovTAvZQLZTWgiW+d2VmeKT
jJR4qGqOMuvV11TlBA8Up6Lh/N0GdNqozzfa7+G9WeffxMQqu84ptuPB21RiFzy0Uevm834Tkrmh
7KXPtW3+4Ag1rSnGgzJmq/Bx7sI3+9XrA/Gf9iz1TE2Bkzuv3jLx7JDmOJ0Ck0fdUGmuI9kK9jy6
4dFwg+ZOpsHuB7mBOGshGsDhQ3no4qSJzV56fB8psnZtXEpESTFZHOtoOPu86KJPScsjVYHmOFqc
KfDxo02JjPjAHtd2FiaD74WHTTnQdmHls2UKIwq8Y0mlskYSlabpwkrOHBZakpGjOGMw0kIBqDMn
Zx0K+C8pX5If2nOOAoTUVvoe6ggu/gNBYU+DoHuS68W7Xf2tBxCY5mRxRFWM8n8t6DgTUYZmVxru
NfrMPZ5Q481y+TKEI/oukXFIaMQW0U1UtmbL1kybhwUDzhQCI85ptcLECZBXHVdxuZoXSifk0DX+
bO/6+pZSj3HfiYOYTIR9T6WAcAM/uo8qdRQB7hKhc+uani50oRa0Th1ebvnU1RF4pldweOJISDUy
XrWvKD9f5uodLyXIxVFzY34mvJB+pt4hpCzNpmbiUP/DmwAzTNFQt2skQV6WZgGYj7p5nXhV10zX
OENL7DEBYt81Ca+WNkpUa4pcvsHBtTvXZ0ppy1CeR160dvy2XFpI9XxSqZ0CHui+7KSN4xYnE8XY
iniKTJf2JYaD6UUevcNQP7NxUMfACJHNf8POvXy6p+yspZHXg0UOuB/elWEd2MEu8gruuCdB/Bg2
Y4GK1Evr4UVabnjvRrRFQVr9ihnrd2N7rC0JW8ABf/v/vws+OBRgG7zgNWDlRiFptizhvW/q68/4
/IbSIuY0k15uzlZOCOqw9ifVXRkzUG94uhOAZ+E6KTjlxYmPNE7my/d6fOOO4JdUB+255+jhfsYL
xxxuf97iRoIkQae1qb/CUckbBwQbqTFaW5/EvaTtZ/Y7OiPKBXQ/i08iDPFIHwcTiVwMZ/0q12HM
QwiqvlO98ZUW6zD01yvsyYEsFnqHjCeIAznwhc0FJLr7X32MhNkC130NL51gb2W0lg2HP2o+lLNW
rmqYMVTD1TIRxxjPpNhuNWMgpP7ftaQUJ6+77qbMvmmFqkJTldXQb/U+Pequ+GwPOfOylMvd6A16
LS+Kgnnx6MeWh3NzV7H4kJ/M+d1h1thfWD7W/J4KxszCd0+kmJKHbyyW/faIewAzTxvrGV/RbdmI
3oRrsWxkTssqwDQ8+iUIO4Ba9YbZXxMwEAIhWnvEOJ2tnI/wUdNFyd+80IwZavANekYvETId8rCQ
ftWg0T3xcN8ampfrt5RFXPr13/KgIV2a0Rdbrn0fRBiHkbTfHYxur/E4q6Hc4Z7Acq7F/y6UJjJO
BRqWhowaKDAcNol/Zx/3zk+p3wWdEGJ7434LYeKcWZXv2u/HDRdc1tD4w1EQmB9kK4VOXaTVv9Bb
z68r1yCQHF9dXe9aGI88AKZf483lVlXGGfCSGCqWtMVKep9J5oN+hQsL4wvKuV71FRzSN+eQq986
eGEDjrn0twkFJxBKT5h9elrp5XMUEhXr0Xexo7bRLviGqgshVhaWb5N/GFvFncUx+W/4ijJd3uyK
q9zoNM/P8KTXbm18i2lxu9rqSY1lvvHl88KPqMEKleWkjd5ytClueomZwTdvto59XbqfoEVqzl4e
U94qI2Y1fhT216hMSxeUd4Ds7Eymx+pz0rbXbS3/57GX9UT7aagTEONa44KrKX+3Kd+opgKpP54m
OTJwLf0KlIu4gMzU5eP//qpY64Wmz9bCPiV4ru/oBf9+/mIrxG/bpLDdxIbmLZ4kKPxx+nAS9R8X
cG4sbq9/2LMWJdvYK9+RBCqZLRJ6DEmGhp+RpHulqVWJZuvo5xwhwAKlEdiViDMMePRICUteSlx3
8/5PO/iOm9xGzbse/UQ9H/l0f//XjMlc5mv7C0HdAqlywjP7Ud1UzLkXp+gXeoE8P85P8PUSYV/x
8mw+f6udFVTSO1jbK6BmFJ/q6Q5Gkfm3XR5Tc61en2Egkvx0Maz3oGMUheJE7z34UxvxhRtaCbJ/
1NCP43Kv8+s7cYf0r+9aZ1k/ZAMlF2czoCCGhsiXceG74gEv5oPtQF5CxY2vg+l/nGrcSBiXlxAl
HyBPbdANQ1RKAP0iwaiXll2W5JQ8kUK/rsSuIl4plp4rnbp5z5/is4hC5d99N3DzCy4PMi4uOB57
Nu0Y39W1uQyP/l0HYgsc1tVv8ukLCFt8lnMIuezZvU77hR+P7IzfCGoPfRapQ5z49M4OXKYxo0ym
gu3i4gacA/5OVBP/hYpecxxIGLFA6J99Qx7dKWCsbz0BUEpoZjuXos9sB4DI5jKg2ybpSI4alUWt
uIONv8bfcuyGM9G2JoFrF/xZIpQBnlGsB445o0NdLdxjOIvZjFJMCjenZ0Qb6eouLFDb7KP5aNUk
KX3DwDAn2fJTyEriiSdwsGK7R5z8Sd8mzZQ64exxLcyPHc581qY46h3DQkzU193DKduOd6SU+8eo
1jMwpais4FongCKyxlY+lji6dy/fq/SxYwGBjPJYbwd8kk+VXMd9EyMw39fjwlthM3YK0TI1ar9G
cDbafkR5m5mqRuvA2mEbgksntineTxx9DZwuQmADhojZRvIwkJN98b/xbdA65iLQcRH4gyr6iHw2
HwONV6F9OkWimv8KufR/3XPImSahqfXhXOguTBEKy/Dp1PofuL6NZRQX9b52TrW/P3ZgajzUqCz9
D9del4IJ+2VGkcQa5hWW6U6ITGGZMkpz1cFhyFdHe1QGfydjh5bLifpQ4fFZJpQYF0/l7OWg8zZo
YYaNsEFKTZk7mOoVWq+YMpbY2HSJcMnC0RC3d+RcRhQlRZUN+Cy9Dmp6oxjuisH9Lo1gz8fqbOI+
0N21kFR26fpjgZ90CsN8b4lowgIL8ktU0KEw+YY2lxv/H00RUZHc59tUOEQfLPJbip9xlhG4aOzH
dqkGWPpChe8a7G8se+Qo2hQxuKjl023Czzg3GFAmXX4RS7124A5IGCHyDFhDLZYnGDNjo2gPfPNv
D+Kglf/t48V56qcWzdz4SzUxmg5Miv5vpLqGKqia1bFRgT5UiIxV73G9KVyJY65108JY62lt2mSH
bnzOnthB8qt6TsMOqNLT3blp1YJ2Q6Agy0NCR3zQ2PSw807iq+AVJbK3lLGlvcH3KE87OHjMmIMq
UPDGZybxepBtA6FLbYLOoI+WZHkeI+bK1T4/TsSScVhQVHfgQ6aeKAB/KI4dQmr7rB+FgmPTfWfX
88fFlUNgRCVFw1V/4U90s2U6/CS7diLbPeJEv1BhjYXXJSGdkWzkpcwJHjUBhY3wIO+loDuf5dzC
TIugHJH/48vBQy/VidSfCnJYpX4OVUTafuFnNGsT/TlwyOuX3Q7kac36BB3QwD8l+kQnxOmis7OS
FqNPlVcSKxSTe3d6XlH+0GDcbvKWmH1W7eejl0k/t22fF+fslSe92TAmTtCS8CeJmHeFwU+S8G2Z
1aP2TJkQLdi3Op3N37zc4jghf32h7Sa0tHDpA4XjnEfqjL5qgWGV5b0lOulMhtPQEgkMmno9XK1T
HeRWMyjR/8OnXzEmfffpgGQuBvOwrQX1hqnvEVGHyGVxgtJ8s5ZnB4fE60OJVxPcqbLyWJRFUscr
+9IG/3VTOFAvS4mTXKnvFd5XStkM04tSEzQIOrWcB/QeuE+VYjuvRdBOlTNzN/l2zlCDpWGRKPLR
x33rNycjekTUyTZV+Q85ZSFbV9pXILhuN5Ev6CfuPj042J6xIbnXZH4Qvxc8pmV/scdH2i1Kv1zK
2xwjAeV73Z3PSTHeDQG//O3HsRihy0tdYvIfGaszX0I72dZadvg6AS40S/CTVzVmtcRLh43jhLf9
E4OUfLGL/pyBs0rLuu+u4bqFVcS01SitFZgiFe5SO+RWEQpgsvErQTsk2QcNxhSh291Uxo1q9V9j
b0o4O+eaxQWBGfThNr5uop020wqFBZpkWz/C1/mO8tnB9wHVpGXEp1knpI2V+VUcMQ5nfA6Hmj7w
SfusY24c/SVjhJGTXAetlMO7baKiZ46a0XHVa5rCIXqbHAGaYsJsBLqv7oTty0oMIUyYju0Ld7IP
DLd3fiUixbZB/690UZUhrGM+6MK/4jQ/Em0dOHlqf/lt0tvjBd6XUcVffzBVx3A3k7rFm4cOzU+1
h6uA+YJNYkG4yjcQqCZMNVxewa86T3cVQ68hsoSfSVUrtueAkglcqekEfC1hS1rj5n0VnYKbOmRr
6LLRQvxWdL2uNnlciWU22yTaxeWbzTMr51msaka+pyjq1QSd4XoZMm7RQvYwixSrp1RoV4oQ0g6g
LBNf0iqNWC1UlyerCoFOXLXeuj53ShOEtgKaCDjtoc0UTLvK+y9k9DVk4X6f5yCbvmJVGc/710o+
J51Vpb8q1bYzwTq7QR8mbIguG8rZSUdCX+E0KaGrcX7w1WjM1loLCD5w5sI89jk5DY+jqyibyAHE
yAtzl0dt3+LGg1lWdo4TMdgUqJcHt6dtsWAmnhgk+9jg1zf9MLnYIodWFAr7XD1qM8gmVFESN+qO
aW9KHnLlg+0LTZIUoSu5TCj9Ahklsz4mMCjZCoqZCgfm4lkuOe7ByWDIHhzV1GfRfVaPbQ/JLs57
BDZKJEBJU8+wFINFGmx/rs6fmDrzHFnn6fg50MQ5lJzLLxQkunOLrluY95flmWo2HR7zxnG3pw+2
DmG/ATUKi1jnVUm8G0mb2369uHMB9xI9xdBKcQie9BXAyC3EN/nlIkszzGunomq7uMviqTfS+2Hw
VjDhb7lBpB5VkjpHu2ZRUlkYUxCDo7cLlPdb2lgyHNJeHNKtw/jhlWYqfIQXj4r+BRflVN0VTnEc
KkAyt2Nkjqa3gKVflohCTUr0NmTs21JhPYxafy86abJo76ta1Rsren6IhheHvjqTzvdRLJ4T5Jzs
+olhNXxZt/5Cp8mOFj57BMWcp8CZ/BhkcDklJciouJ+cbzcxHepSrtPoUlfSX75OGyaa58rAq/yD
dmi6eStaRV/A/STZ7FfTwaqX9xY7DevFifGKE5WZG7Dqowb7fpODc0UpxN+F/mofOC/TLIl1B12s
oytU8mwNbtAWke4aPMx7jTIVC4N49jiKR6yZvuuRiJqAC8hmxlcGHV1MV7TIoE/ni7COjC8/8gPE
UfkQQQRUcaa1LIzVW4eo+IFf4xYW6xN3Jv3t6MPP/7VAmfdgxfq7AyeZKhVarvoN+xRQv/W88Fas
fC0BqI2XU55sq2FCWHII5rJjXZmvldPIVL3923SDYOVJfXVSyp/jSR+zvHfUHWV2OQfpwLFA6y0X
2rziLTJZQipuVrOhjrPBRMZlblwAhLidBzBIb8Bl7UmWtIIG8M2woBKYbg+gVTOUNXGIw6p8IOyH
4n0BoiySkRS24hC+Hr02bjFjtQWIFkVbtYVMwWrNERuzm4EwRmnCMj4EKPcpaRNDLLsFDI6IQpyn
sTCCuUWXZ3SLtni1x4DK8l6IyV4+VO5vHyYCLb5Ku6RZqkui+eo6zOyifY03u0oenfydxQ3shQxo
RKmYROj5Eedu1izxqNSQ4Al+9yOAfJ0X00jQPkneZc0fjFMi9ULV2/gk8DeXmvY1ObDWdaA1EzSz
b5kRfdGxUAcZxeN3hKom10w1kzzrm0/18nyqhw+jGe45lAxuxXy9YRUoDlmZpThEP8BS1hRogvq+
IW7H+CJe76QeLbfP+NpFjfPZ/K1O+fmmSZlCGIGvmPLyFA5SKox5/Ta3X1+UFANsfSIAHa+74q7+
GRcgt4T+bUup0ZCBBVEQ9Qd2YAVzIitG+c58sJYFW0p7uPrkorl2N2znGXrCoQQD+pogGCl/yzg2
4yKqZzanvNHH0kVpJVYTmTgFEJIrdEDhMkdVJ8fi9/rIU5CmuvuUw72iZBWaBibVA2T5kEs0n3my
lzlBeQpuWm6LZboLffthTY9oaDoeCNfpVl38mltGQhz4n0GUrNqV2hhqiiNb8gXXztcizdG9+KD+
8tPwuJjPcpd21sLLiUgjeOf7n32Rh+VbUc99XzoEWLwOD9NfLXzic4TKzc1vpeLdLxoIu98Ti5cs
V+kKAeR5nEeVakvev/8ZG3HPgFqS/V4jN7BcWXdH9gNnnjBuvAWkaCaUq1DidNrVh007T4kG8vvU
ef8vq7Tcxfvc7mh3rJXk+NzHmwROJGAj1PxY2Sy4sw4nMvHBWtFbYVPNQbkRFRjc+9Q6k6Hjr1jj
lbINvXK4L+t/y4I6IZ25ghJELc60dgqJPt2c5Q4IKN8K//rOT0XOjc2ptnZD2Uid+FQUI9Dnljw0
daCt0PtV/kozlTJKySoNrn7ZgIj2HGwLfhgpHE8mHVnNk/PoLNhurLrj4fDh4YY0Leo0GAhaqHFl
VD3Lxdoo2NUc6Lep7GDR25vMy0oYBveCEjWRUZ2iwth8i/gSHhpxjS1s7t8zebK/rvlgdjfEnAB+
cF6WFB8ExGTEAwdkza8ITmF9kNSqXleqGlJGajzPzFfOX+2plnDgwQzBg3SZAG2cIkDyNWtOLCFG
FmIPwdcUVA9INAqm7L5nka1eOeOU0nd0tpOofQaOl9c1Dn330lVLU2dNKw95azFByfzB5GZn9LyJ
ydN5iWAaaqNZcBuwoMVua+rDjejr3M3HiTBTQbcl49XWNVzcukvU60sqYFtabYAP2Mm6KYRPkx02
1wqU3xwkrkc0eN8PJVmcggQdhNNXwn2gpFUUbwIvbjTSc1VBn59i5VEx9kCpMh8YoSWf9NxMl5ZW
jMssQOYKU38OM7FWBrgp03TrDPIKJSwJoRbf5WraBD1BlieEyojcLu6kOHgKgA2fIG9S71GodEth
LhgYltyzGOzaDcCLcWA/5CICF7/mwEbhxOx5wVGgBvQWJsrIibcqbWoGjBMw/25bDeL8d+8nRGry
DPq87WfTb0nX1yYZ7VSWrxJelX6tO8bHiYatdLykKuxx/QRj8/s1T/Fi/GfkcLu9lOH042RexVqE
04aTem17idLTAxsrB8CKy/KVDulo3YwWdY97oiMIH0AcqJVVu4PGQ/nPF5ynVcXFOK9Mb9+oWHJU
iMevvLlAbG1DG6r9cJSUiK1yXbDR3u2ViPqyw/YfMicJFz6uuZX0JjUWfr99L1Mn4nl/9/eY+p2t
xJhI+63lBGblGWKfosGfbyx1Ad6wIuN4eA86B8VISGPdOQaC9iiS2x1tkwtGX+HG+Oj2xFhmMbWu
H5fAOwM5gyxwBbqVuU8J6OXIl4nsvxZ+MRYFcNz9UhrVB1xmgheQwTVU4nYQLR3rgrBvZZnJKfLO
Q9Fgbgenzni1ToLQvIi7+RlxReitPorMWxOyqxhvfCKkn1I0Xluitgi3nTdOiPwVs8JEmHvfPiO/
sRXvLlObE1U1dn3j90XZPTiAtPYBmG2ADyBRPhzxg0JXMtpEVwxxpCnw57ce5RKQww49+8QyuxZ0
ioJQfJWd0Stj/we1iFz+yzTahwm7otgSFtPi+VWFeyVsb+j3GoRu7ZTjYFQlGRK5dpv66ecCAIxG
lPw/bxlwhpBF5X54Al33Rjk5A4tiTM7HcuFuThpS/2w4wT/1tUkLDuWLIGyNODZbPF7H5i7HPo5E
KCETQvQdJlF63Ub7nD4QaXMgygHBRj5gceWg+Q7GrZjRLzPtUmbqjZ0qw96Y6dNDe7Q7sKBbNSD1
EV+Ui+vwVpIyZy3h0f1niI+rnCdR/zezPUsG3pM5Ww7RaWWMueGgysfXid85xbg5if4hBbtsEsgL
WceLuV8+csqrKHq0q5ogujocG1Uo00zNXtCh0RZ9I5YjywKTbvE0OUGxERXoFIUmT2Uqusz7fYHx
mBJsR8OH5HbtVHxAfaBJBSdjYr1YjixIGygfG3vUasGX1hon15o3Wy63IQfukie3bk//08C4wiwc
19MQCS8TSL6DTFc04cDW3DgtVy5J3GGdNn5IltV3j4NstPQbFSRgRIWJa6oWMaKIE3QtJnhWTXFr
IA23kSxGdn00G3bOmku64LM3ez+hp/slw5BfbMYqTMHAVc05S1cL+irpzdtHx4pi222lbD+T5Y5P
5sBwSF2iaeKqPTSICTc3aMd6wirfM77cX2bKGVv7wrBxcBehkeK71EMc1Yz1qsodFhkU4k8zrf4N
rgi+0BPJGEblRGcNwF0Ogl3N2tKx1T2J7uqSEjmivTWyxobVSoQkXQ2ooYv5FqdzZ3aJA/4g8wfD
o3R98JGhHxbUmfDU1e+8IJaQUSMwrcz6UrNN+fvQPsFkEDOLv9Tygpm6+0ZpkVrK3o1jSdR5O3mp
fcjexp7ndMwnZY7YDsBR8P/t+VAUhQAQYCwNjPu3lkKMSH8FdZYxZFqrzjLIGM1AwMciLATZRjlk
pD94TlZ4FIrSJwFrqyW0vpE0mTz0V7xS1NMFhnjXuakFVJAVZjNT2UFBTqi6SBoHsNKI7zFrEOi5
vnA17pqHmZvg2mGE/tCpUG3UwnwU+/xhSMsA91rDIQqrJdX8ibTnX+59+i6hPEuJf3ccuh70RCan
zUKlzJOgXegvW02FCJ6WcTSxWbydFIM0BeQiF+xrSU4fhxtKKKHmhjXRkwJuBScKWf/5N+UvICSu
d8XSfehfLzDnuXSNZoiQqjmE4FZscH510Lj4xGrWyzUxEKfJy11I3a2DAxfFHLOnFM9gu/sVNb9l
R7zXLFu92QSjIvnvmNQYk63V5kvNWXRvPIW+hGJdGuXco7PaNWC2s1gzPFJexND/pTmcvHhJAkHJ
2scrt7i3UEtr8tdOR9buLU/3fcJrTbavEmm/Gf2ckq9/l6dmdsWaFruAgs/by8dUwM0UukBVFGto
g8Uiocf05n7rIZ6U3lsXj9rjDODD8uzPumutpwoCMCv5jX0SdrPIGYw2IdID1trbMLevNrs5LSoz
90EIrL66eGfBlECbNyi+mm1BhW5ztBbMuG4pqsDEm7l/lo949uzPT0ttmIFhGi57uXoYg+iF4QIF
6AkLirrCXzBmcn1Sl79ufgJJbgElQq0PrqTV/fl/vT9SofJs6amdGLQrYN5yeMEu7uWTum7YO46b
UW5drJgmU7CiE/08OMZNlLHLoZqZJgOM53Q3qhX9dG1bSblCASqE2+D6VVLHXYLse4dzAvC1PqRH
fageIb5MzNiKrFL/7/E/vnkI27C8LD7x1GwfbMlsLkRCsHelS0fJaJexBsZfOExQ+AqJ8uZksmTp
n3x8HpPeQNXe/0KyTmt+iAh8//KRPSk45idTGoXtFLCEDewpa8pw8mkuHKP9yky/o2v2xMXEhgzm
P/qjG6sPoDtco/flFKCF7axG2PY+6fSkLEe3OGc/QGlK170s+9JAoJQoy7zbsIBe7MaTHieiiyn+
buNehBNp2JPMi+AtmQZzBVONhJdz83EksXM6oAlqxDb5GEarL2+ZFBXoayP7Aqc864nCuEJRaRqq
So9hEbGNa9ot9vFkdOEoPdUe6DHO0gc1M+EAIQ8TrTswlONcWgShcULX9KyrHQAg80A6W3IMaFGL
RJDozGMJ4hY1h4fX0Ll8taj4UCnZg3nGdRTIKpbwAzesGaETS8OcDt7uMxj/2O9R4UhrClFhUAJn
Qlp/BVjrOHvSf5Z24J4ODNxS6hu71dg+M+HoVzjJE6Fgx8NNBMV0jSMB66iJTSqw4qe9gIJk2ZDu
XDpJRIMjg087c7BXe1S2ylNF2bpTs4SIYvboSeRzYpdPeoDLY431oAjI2IiCjFxiqwYaZ9v/N5wn
hURuvD5C5yldpQEDjvTveg/TeXD4P2kzwx67gpkBzeN2Sv4Puymf5RUC0vEHxfOh3c1KWQ8lXmxf
ccS8xvodDDNCGQfn667PD9RPRCWrOm2ClyxwaXGhaCqCo0q5kZ07bRwS2u/XomYR0qbJ/OUgUfXy
0JY9G+vjfTXS5DgrK5+Iea1YZBiixp37tKl3HRu2rhoAR5talKzOiH1sDxdOgJwBzv07ht3WTSqb
Z8G2/2asrw7Q1+Vtuz3cc8tPeFVOABV0n9QRLATfFXV02dmI5efSIPTcJs3AykiyvkiYMi38CT9M
pWvcJTTCZarluMijVsnJi5rwtiBSytQLBfO2PbL02x3o4I7g2AevKDhrABLj0qcALrB0/We0G+4q
KpwVOdBxYXILd+dN6zC2gR1zcsTEGkFIq43xcTBziE/NSoFiIc7euTnTDxewHh8w97fNNXd3Cdsb
bpEwpDUXARfx/5QNL6b2WMeEUugjoT8lj9NlktzhGLNzNz+rSVL44yA7O1wh1XCvGgMM7ujEj/Yo
SS2K7pEpzcxYgMl5BPW35Dmcdu9WWEfD5sN60Uma30UUTnDJXioq0OlUY6U9PhvPXoYltWxCUvIb
b6TJJ2IQdsqzBepKjfy3qGm3MoE1MFlftTWeynpaRLmqNOXV7vz2c/LFG/y8qjz4pnvqjDdRiUF3
sCGCW1z7kWVeL7Ls0ta08/T+ybVWHd9VfUIpUFy0iW1tZNYZTutWrgpg/+CfHwcyKVXGx3gBzbQt
DLMPzV30P5KkoW986LUlmc5xOVz4Y9gZs7YKJIeZpGn/lcHK0KVfJLvWsdGWTRlze0CJ01bjdNCK
7uXAbFCAeFqtbP/0KbcL2UIvmDjPIZcFZsbqjvz7+AngPT+Lx5jBJ4WTvAuwb9jWVbhvgdG/VzNq
nxST0Q5NPiXIDLdHZUhs7c3LLkq8CZr5+u8Sru7EAV7bZ0a8tlv7s7xJNU3hnlNLm3Zz59lu3Drk
pW43PqYZthJbNPJiL960AZ32lD6eVKnTQMlTcRAPIqBrt7DZEwt8gF6uizb3HCr25DEHfO7+0oj+
7ygmwKkAYEeJL0ch67phIqnQ2dtzJGZabeZX42YWCp8MCdJqZHWmtoOipmK8j7e+ECfh5jz4rgO+
H9QKM3RywYXi66xwwmo2NRLMgMlQBvdAz1gCVWx2vj8SPHvWoNDPJq08oyc1rZD+JEU/coDmoBJL
NBmiV8coSu90qT3/n6NXWTvDWl41pY142X4YiGNimCmNRTz0Ss9xHir2jMK6qQg485c3mAkfiTWx
Zdw5YDlw+n5eZ4EYcNwYirvwPAD20mmiUs1Av6+hkkll2qluJ44kEeSYzMNuXjD/ldcqD4yEgwXO
wOscTMxq1OXsieCB82mrQ9PYGI89Eq9e6mCOBaO4jjXXuXwo24IpX8iD2jIaDhyXYk+hYblqLxs1
cGWHiqVtHNIbEqGJGikP9s1T6PLU7WaUHP8rdTBY+xHIwiZ6FdNLUf094rSkKeGitffVeAkl5dmA
QIlIuQHlJxy4NvsGx7I13YN2nXKOTi+6EmmBwi22RYrtyjr5IJNnuDuwcToYjmzv9rRkSUACNjcQ
XpMbHNf6AKxNN7eAUdBKByOMeC+4iSIb99DNsGSYstx2Vo5rJl7LHoHlL8g/3lmB/HJjrPtoQg53
KHE643jqjFpv+0V86U03cQGBtufy9GqLVs4gSUR18d4Q6cjNq6ZQxfuD/VDPpH4J3dh4vZvDZqvU
1TzFiSgrFymcg1XCQ9YD5grZ5u73tX0XWVyYXLO8XA9hspHNrM/mSOwv6WiijJiqAxJK3gh2/nrv
Z/FXDFPtDo8MZx8kW3SRgDrL82bUxLO8iOXHBC6z8COY65FGRjqXSZG347QJRRJiw3CZCJG7JYc5
bxncNsTMJ66UGkIrXHJXfV84Zeo4YEwFT4s9DyLFgXHxvxdh5r6p1AwDJ6/kWOrdOfM59U38/2Jk
xCKcABs2qJDIZk9/pgubC+7B/cquUu12H55N5qDs6SzJHyf8s8T4cc53o7GkY8crUvGWhxyasjdT
fH32DNAT0N4TMbLQjZbL7SFHEQ1vDKVtwJlT1QaoPlbrN1KJ+3T3ebV4zQxSh82hcnWvEfLHgqt5
hob0/EKFcAodbkd7fVmWW1KJVzUPw70aaWZ+nPHfDr1Msya2oRjOud+R2ZPgKp/rej50ChCxNc1T
5FjgmgVnBnMvVvyH4ZSmW9UABSfqDSPqLrW3zCA+PA0EoxN3QGqIBwb+v5Mct+bt52mz41ZCBycU
wlEYpSCAaObacGo5z3XjFoNYfsk82DAGGKqsSSR2ANXcW5Ac0IkrQu2bUGjF0C8eZfvTUnj7sUep
dQmf1uDtXSlN2K7rjNCH4JK9DpFF5R2scjfSTtctcRkC7z5JxwILX4MRmrofVzuHhtZq66PnrVfF
jS8OJ7iyRLCKoyhvMfBzK6KPlH+WAYUfwbJcqgZ2xC+vcWKD1aP9/Lc3CyvcrMr8UmJIYQA1Om3Z
cATWygJ9FXy/R/KCwcmZRWdrYCmpZKSzU/LZJNvHlaxkQqDI/Ky9oX6XixlD/Bd0SrEscVXdSiyQ
7IcdYPvIbq4wlpgHrkehmtzIF+DNe7Rj/YgbH/PN1Ig/P0VjsXR5PQux1u8b58bBc0BZMTh/4Awk
FoC1+ktoy3/lLdoI+/uPPWgPmu9N8Tg1I1TAVGTlxc5YNj0CaAZvtA/4c4b9ZAfPPaQ35h/uJAzA
5ODTCN5NlQiToipCNI/VcCGOxqr6VLsAO/f78Vtg5G2YiZ+dXocYNZUaYSGr0A+j0SFF7GFeGKC8
txgyRv+jQlLAYDRwnKI70sfDLMhkSrXIUKDl4gOOolz33WF9kvojpxGHOSEdaQzIxbbywSA+IbZq
3T94jpoMXN/NJoO5GvMueat/hx+W+L877nUqE4z8fxucd+wEQ9gsk1KUOhARo5R5RaBiCP/Aoyqx
olDdn1GAW40pKf6JhuY6Hn8OA2e2nr11l167SihWHkIIk0IsLvJUSMD4UpF6nrujrxc2Vox7P3zx
xwNumF2w0y2kGiHK5tTaFNXxGRulwMuiAvkXnv4ScGbZtF7LaCYzxgkBj5a62XQhP3IIGok8E24L
g+7955RG/DaUi/VH+6rJDp06foDsILjDp4hPQ0MsTsFaWKh0WgDtyqoBP7h6kSetH10fBA8jKMA4
gp1CPvDi3qGwx6Ohn+965Stxt4BxPxF/DHwZWU8Yh4FQdFHJTecqN9xFyn+4NkuFoknhDqnqNMgX
kuNlSlJ5hep0EuTfqUFvlYi7xwLtUh7OCYfDNhoHiQuJaDIC/2cPwBwfE48CC1OGspR3rIqO8k0l
tKxsNAVp08zAYP1a5n9pt5Ks8qf3BbGciylVCFJdLusXtZTjpI2dVyc3CIX99HulTvGEhYVvuU90
JlOc+ZZDeD4iwkLS9zWLco8vtnmLUMs/ee7+76UUYaJsc1n8iPVUvXmx3WhAYZ9g1NQetQZzP6xq
+dcGW+2EhD4tUW4W43McQhdUI093iDyS1WKeCAcCSbAQGlaMPOA1y0D3VKCwVnhQO9RIUeCYs+i/
YQE72UpOQYhwOme0doP7oLR8Maj1UOWzJacvq+98xgFI42aDKupaNXkVD5oun61m27i9NImxGIzW
zdlHZTKGv27iZwBsW/f733eCJbKZniRa6Cm/o3njH6kEozUEjxN0lDFdSHxZyIQs7Kl95bPlYxTu
ZfFpdR85hiVMpDvAvY/Yhw968VJeUm0TxKRxNvMUwg6D/9imSsItuYg2di317gm0A8RpgTnjN65O
rB2/wPlgt970VgTGKz50umy7JPfsOppEVhYGxcPcy87tABHbyny1u+wEsgFHCl14xJ82lxykF5Sv
X1v/dqXAsDYo8eAQdyw2tP4VMIvjmBPd7oVjrumkzsfdAZCQorp9IZra0xa3V55Sn3IbDLikdsC3
aLtrGCuBL/VQLyAaSNYSsJuzzVA3TGR3g0x9fh1QMXiNdpa1L7FAfX3TO7hgXDeUhFes9neF5oT2
uIYajlsuTqC8famOwlE4z4kOKE+M0SYnIQsb+6uRUmyToM6UX52E8ajt+ENrpiFvuBlvf+FWFwtf
TnJQ5Wwo24ZAVfCj4gV9O6mcn7sqJYWjm0dhngE2RSmx6aIzmQyn+W5f6lVZNn2qAFr11DpUW9n8
ldU2MJHx3prVms0yub2p6qfBtJ67+GW81Kg96Uarr/ks8rvPlwFbBLzC1kn9Q34yy82Z+romMQwe
uq2WCeLzLTUaZ8DvFoqMbS6BeUh1iGqKOBcLHY6z9WAxL/DMIHgvqpWMHYauMDWeEe+majVrGInw
bFxBXyLI1WGQggqeV2kW8RKXToxm1q8kL+t7RD4BrQzC/lWEa5FH6pnjNAiILxvqSYUdJut8Le0O
w3Mr5up6/4bcZdxygKaWw9fW/McKm0fTchRaiYlsQhE62u6sbuR/1vMQRizJar3pgLqAniLIsGsP
jyRD2QsQ5usnTJ+3RbnSSUu1lgVpFs09lwe8WvsJTi5f1FUb4mNvapSMOgscXOGiR3EiwWxPHjC9
YBaeqXuHbR8NiL7m8/Wpdok9hywJ+5qhu9NFLmGlyNBVhGUXB+AvWR7+XE+bWgdiQ7o6pqvB3Vi5
fUb4kqODosdpyAH0S+24dcNmJIS1tE6mcUOtVNl3nRwLsFZfApum8hksPxTgmUQozidQVlr0nRXC
IRxRqATnq5mucFBOKICDGX8zw2N3aItBP7Bq51mgm1hdMe2IPUXh8AcxzKSlvPpRTgdPl38B5nEo
9GvtHHLDixzi1PKNTkTnlgxxCxjkDOEQ/4HxJkod9NvQS+C3M5NrLMKmhQq5mkAHAoKd7QimEZCX
vNh//WeVFsearzmmmfJF/Ur7jWMKbJFPPElG2fnFgFFb7pK5mR9w1TO+MMoIIxIYXhLhjjkuNjz6
IjgfQWvnjNqN1kORZlpN65REKFoRHdpVSPezqwksfWopmkDQn+F7tNxBS4cl82SlNkpZX1CL+NUe
iBZ6nO7fCQ8RF5yhuOmCTZcGitL4hZPDiYuI48jXUSG5ep4Uj35ixfeHTIQTDVwV9raBNnyRo58S
zlsexxiVK+M3C6opJIRTl52eo6BNCZKbe8Ndi7pVO/Dq2FpzsMURlFwMu/BTaKjzxjBdgp2fLa1o
lxutqqzEpfD0GN3TBgLjqdCTZV3y1nPE6gn/A1h+UpfLZB69GC8fBcWyaP2itAWVvHrC/K/LF86H
sT/VXqU2ppeLuWoNrNm7lIYctKmK4+J6nkUlDy3b8iQFRQlOiJJWWEEtlg4Ve0tzE2ykibTJZ2hx
RRCzHXIp6fKdmPvRVcRU6242GdYAbraP94/vbyESsHR+Gu2Z0K5ZW6qIrs1cZaHYcC44pSOJD3d4
cBF3VWSLNb9m1fB0BPBanrgutHinfNVKA4EaA0c8Nu+6yl4m4YirkPCAbUhyGTPXqxXsaIg/G94d
wSuPEYRbSznX6xiWGN3PPzQbL5mSAjKLq1w2lre5IUJPr6F09x+J3O3XXK9rKSt8u7pyO9vppVCa
qJVEXBayqYRIRlmrFsHN+ZZsN9KQ5vcvCZwPyA4YIJuijH7dp+Gj1R2RgE04zw7CQ1Z5BJqaX4WY
Q3CKHHqiGouoZwt7P45oJD+1aryngPWy7NxIDt5qvKwUl8pWNGiUL9Pj7QdBX4IHM9aDXztXYXD0
yOlGryoKk0WsnlXlmCBbhap9Wz6UrT8P70FwWb/GixBT0TqjRWh3Gshv+TCPTaJbwfxUsBeXCYPH
x9mn3A0nftVgqaRtDalVzyUdH+WBALtQIG8TUYVD8ORKqIHdrj5m1mbpC62iwkLF35M97sN5l+3o
xkJbhbCOjW5ydHMsiOwJVKq0DsPVJahbViynj5mbz3Kuaugew63LtAQCUI9/fNxg5d9iFA1Z9+EX
5h51KwaX5h+fiL7UcopE656X+KgOdKXOc77/EiDVcP336BwWaGmgtm4oJiivqXDhlNKd8Shegswm
jle6KVY09wNq2pllrDdL9R8zhfGR1xnyFUj9783erdpdh5u6mTschm2xXH1ncpGiN15zpbrQXLMu
xOLiTVLgVT8Twwqp3rrV70nWw1lR6ZqIoIRuxUsmqoW1S6z2nFOXU7uOImJmmlSNufQTIahk2ahQ
9uy2+aUp+Glguo9tkrI8Wc3oSEDvTUY8hVQXmrp2WCRbJwg4b6wSQi+AMpIFxLhnPkPuiFgn0+z4
yQo0g1crkeN+DUOJAXAQde+PqA7zO68tIC48J9iCnozdZsU6KyE/UrPhCQK0H86ECu51p09KAR1t
8yYMMXqMoJoakDsMQPBquslsmbIvp7aSwonaqynQr0pMJ+HZACQjznPGdP1yTYvQ7ucGJ9P5NDDm
r+Fx9QYyPlwCy9zdwUJYTqKFYMuYBZCrpNXuIN3rGZ1FzxAgc1ljdspjyq3edbnk6jnb/YAVy335
LpOiFc/Gm9WwVtfD2sbtRwtQuAnvQOtmME1MsKhqFANOQqytiBTIyywH8rl9YOG+DNbsMVeyFuKR
SyiBA6dXUVjYpUK/JaBVOhjRM4OxxFd+VAYNi5zMULJlFZi4+G5SWIV4K1c7Xk7Pk2D+ZxDW4HVW
OVcyeQeGUGJXHZNg2M9bYVd3kYoAQpAnWUXcuTYDUqtKc359rrfBUQCuZCr1Xn3lggMmC7QmHa3m
eFmABoJWWDRY0nMyr06onM84JnVgzZZjdj6hoEL9koeE1225um7Uq/kjD6NcPbtV1PIhJdVniZzt
/rNsmn+ZZqMQjtE8jCwmxBskPOwjYXb6qfhTichhGBdVYhaYDPKX796Z8dbt07jOtcu1lotwM8hd
LbErALRpDrYaJRiW3HGfFQ96BSOqCjePeXvl76oOjd6xr9IKkGfGvNlW97yeEGoHDs5Y728Fq3Ym
5PFCJN5BWBpR9Y1RLriG8jEOD0KyzOcaXNTPvDLXQLFogYK4Q3SBCyWBWLUt+RxZctv9dOjhyrp5
Fzz4X/4oT03ycJm7e0H+y5YlTtoLWg+I32xyIUueM+3HiaSwchYVcpg5HaEDNFtXr8/9eXrkQphD
O5TmJBYbj3QGQUgP8Mj1Cd8TjyjnMGP9jXO3AMTGDBp/0Des4VQnBU4KIATJMlcCQBLQYWMQrgcd
zmUD3RyOhjRTxTLY4Wi8JQnGzVZz2GoRz5YweKjKGcZ6z0ODSb3I53kTNnhzfGqaVP05nLd268ca
BIlm98kbeGrs7r6CvUNxHp4kkU7PPxePBHnTgGcNcKHCAX2YZSDpvvBX0Nx0hbNqILoq4vDBVF01
ezdfNgyMMtYX8jelcmSkJISTSL+f4//xBmqeg6TpBJNgenFjzFfLVqFcsckAz0MJGTJWFhaR1wgF
0XLKzv23oM1t+tDP/mRbzUfgAfvWrMUHV5YvQkPF0JTGyBs0PtAtulLM3UOgdn4GU5KXmffsdEmn
1MhE0oy2fJc7Oc90ShA50HJQB99u7pJTCBtjsOMnFvCw2lIsvhs9+NFgnxA8KTdtavJkCnP55N8g
IADJ+E7TIRk1INwwIo0kxuD5kI7jUTBSiCDOcfBATE04qPhWDm6fykqlUqm0iIXJymVoC6YE5gRI
LcCshkv0bePL/d8DIjErKyjkTZtjLGRRfDyP6HDo67i0EFMc6VhI24xzgEaQDTM42nUk7shESWZh
T2fKjhcSoskzLNJk86QUVxnPLggp8rdsHf7CMejT3HckrIlcdZZ2zeAgEUetGlKspwQCy6scGyJs
xHlPfFv1jPi+UW3b888ss3vwQfu1X25HNrZ3cuS3SaklC9Tv1hX4hjcTzvPbrKG2kSEX9kxqi2Ha
2x6PhFpGXLrcGmZGEUM1s3T8FUik4tCeeBGRpxahJR+yOn1A+hvv6XnOf1z5s2meYnQDaad1twy/
uwCW7s/InMP8gVMW9BJcxyCXnIE0AAcrpjiAZD640GkVTvtqb6h78mb7JM9tothPy/qauRujdEZf
Vw50cWvi/LHpSTlH3dYtBI9gGy/IYNmg00L8JF8FpHyPtckyeqzJ5LH80zEDcQFJTg+ttVheLK6a
PDHO98qsokJJqf++3liup1KavYUvYNvjhTHddZ7O3OPWh6lz7qe3sU63iqapGjC/CbfU1O16xG6U
Y4sE++3OBuN/oV8Uj1QUIqE3P6BtKCkaSrZFDLCUd1bO84g1zTwf2AuNwNQ880dbIBAQxmqi8Y/L
ywPMFEtC79HZ94QLaIPf2rIo2BZxbwE1aGZ8dc5V6xhIam5cVJJA5SUDHOBQv7uEpiH6iJKYhvnw
HqXUsOImFeEH07TvylK05/dn853LDpZNfsV6+9uAd2ALsjsc72pO0VOw0bXq/1lJZVAFgXeVZOB5
A9JWp2z8ZwogwsDT3bFVO+Vvn5yl7Td2VBWCR8oRSAKAFLmD2/aUcR6NwKIMRS8x+CnBgs+SaQKK
13DbQi/0Lvn7Ti5DKMeTtdW3lbLaf0DMFNmfLM/38eYXoVkE+B3p6XihAkuF1sx0OZ6d/NyJl7W1
xIQ5f5VBJgZ20vGHEyQZaFqkvSlB5x39qezGAenlX8nCenu36+xcsh7ZE1Ve1AsgSbafTAqKFuXL
BkIGvdKxb78nuFVIkptIlxnAhGwd7noK/Nb0f6bqUH5Bk0lIHLtAYP6ksUpt80TCei4wyelYY9jX
cFgDCO1RihYgRF2Ay+3y/WcHVReQvE94dPXpTYzx2qO+gGvkwo+LgP19L77d/tva/TlKTjH86jbb
7sOe71YNTjvRB/qlK0USJNpDL0gYB/CY70z+7x1CkXmQ+3pBFRKntBNLxqvTw0859mwUE8lfx409
+Tg7zgcfjpg5NBhS/21XJS5hfIQgsBgZtYEs7ulOGNHImgVqk6hlIIxOlu14JZmWlGUSykIQB11L
lkfJLESPheE2T/NvlR0BZ4+nh71TnneBhYUHnrR6mRr28tChZJpivALIxi1GxHg8NOXCMTq8iWzz
azAP2YuslKbzmUWbDjzDd/SdN8XR6TpmuXAURJ9zuOPBh+ptZx7ZTwjT0PTOjgsRXuZxm//cse/d
JTluTkNPl5BVbCdk9hg4VnfuuCPafLRZN3UwUo+l90lwqjH07TOww2keNSKv97dVrg6n9+Tid/vt
sE9eEsQ/1EeCXBKU0JO7CWC8ZcYVOIUDGIEWbiEMSWSHfeyGhP17E+DHXGnEYgBF1IjVpEH4zIHn
o0jLd2hVUiCrDyZCc7FCafNOI2Zt8fW6nV/JW0HaNZcYCFKqeRUCvrp/nORnKoaZVL7slG4uXham
TrjaZOOZkwa0MCGZsZcxb0VQRbX2SzH6ZEX53MuNldzLOdLisZwrr20pkiSOD3DfmB0+C7JlpRoQ
PcAnl2xKlEqyr+cZBaGKHJ4VepVXrgyBzhQhQPF7WUlZVtjxOAzPYXEaoOC/695irw2aEXcv99YI
bdL2b9RrPgqczhAj3hohDDotKVSfsAXbn4XmuaelwHR/RsIJHN+WTSKfjqVr/pTcyTn0gAhCjO7C
Xiulufq41gmpto1DJwC3uisSp7FSz7J5qBodwI1QqL0ad1r9izmM+JclE85+t2LTXjWQjXv6Flzh
qdBrzy/fRCh0nRXkcc67VseC7et7PuXO4JKYKN2UMYDyTg4D5bx5/Mr4yuTlzD3UMa77PWO14ium
oN5U9MGq6wbXBKBG+DHVSkOGqdi6tpUJRDMcm/gHF67TrosHCQHUp1audDAEFSq7d9966SS1igYk
W47tnIPWPt2aL1aHOf4vJ/wVeds/VzWFoY3iJMI/JN0orPUQ1aVDUVPU8SCLAYD4KjXdRwp41YUB
Kb8+2sVsrO9EMSQnTXDvuPOQ+uxNYnbn/OGFY/Xo6ETDCb56/SOBrWHN7Kn8EyfD8nhqEbA+DIn4
vN1wI5BnmvWKMw/rioLZQpZMFCNGwLNBF1zecJQJH/lAxwqjTxkurlPABdiNN9ID+f9Fsh3zpqln
ejJMXN0aMlxWx638sbGUU2RPUdT7s9J7wdo5QIVDFhle5pQnNI2o1W2jiukrk6+AEFRyxmw1ojJ/
FZ/w6bV6GaVAczzcN18LALMpZE8o5tX24cqkFI3P650XsanAyd0XJzZ7QJ6P+BE5oKyF+eesJtxN
Jd9bKjxPJtUbbU/JVORd3IcOWW2MIYIpr+w8CsLpLr5ZssPuTdierIqw9lbKTR9BA1hHkb8OLic+
YMu3X7BxlCZkqeusobKDW3pPBSA26Kv/gPLeZ7585vvKH3HqrW6JwxYwtCSNRo0iOybcjkkOl7Rs
EaBq45jpmSYL5Soodv3NTE3DH8kF1THTxfGBGbqyvYESQe3r/wTYiWFnQyuWdNDtOc6GlFQ2uTlc
TU7q8+0H2B7KyCs8obmOQp6uGDL9hAuQLoid7wYXpUoAhv/VinsxGc9qcJMd3zWQevPRmr/R5mVt
2ryc1s+jsGWniIn7NiiET1YphWvyOM8cnizerywqhSl756MJk99X/015WbBRzBC4HZRX0HQIEYbj
DTwaKihVJFnsVg+atsE8gVz7W/z85F2y9e//89L20SOygovHvhBSeuF8mWhcKvylo0Ic/0w9709I
rYn/Q9fUb9uP96whcpY84osmSa3UDNPZ6CwXfu6Ynojw3e8aHdFbS2U1cs5tmCYeNGeVZ6w1c1uG
76k60v+YomGaRoBDfgwMxt1DjdCVl48pRpGXyUYCP9dLC7rrRxZfoWYbPmxLZ3tkNfIgcOGGQxRx
6yI9siNGAe/e49uCTxdBlrS/kaxX10t6LnP6C5mCnpffzAqGSlPd1bxgjff+BMRVbdq0iJRu2hQ+
Dn5MEsiEKoc7viBWBFjG87ffueC4x5SVcsTQbuNrMutbKVovywNIWWJooB42gBttrxCCw/5ytAVT
pOWzP08cLGfxYtYHczYF4Gtu8YevyFfb/H9m7zYhNkt5bhx9dIyNc1Hd49QhVulo9pZNkuRnSFHT
TDQEkgwKO2wK4upiYJndfcoyZN0m6nmhDADp5JpEdGeGe3Q3ujFDPjE8JQhCkIdFodPjBIP/OC+u
p57eyPi2mgwgcr12jVDhDqJaJJmpEHDDjSUxieIrjYIRXR8aDIUy1Dcns1CTaKtgjoJfr28v+EBZ
g+b4WXBhKF6PU7ox6wvgyQAgv+YncCmsvs37VeJAO6u0lFT1GRBW/knKSmWl3nhYqI44VJEEbBXd
jHtxaGAZXyeTVZdePWas3fQRRWMEFPP+XlA5HFpiOHaeunr/VatGDNUcPqrylM9uGMt54tYWzIGf
0xg0QETwgQ/fmM35RYeeeH6FYSDXKqlbwHcknrMNlu6K0kC4yfLk+rpn0dp3pgqAJjJH4ZpBr1i4
KsDQHGU6XOzjwkIuccxZ8fLObooRhmJ/tLQfRVxSOPW3WQ2kWUOvGy7nGoChk12FapIttufa3xs/
SqcSCGquqvkISvwAr7tZ7LjxN/G2PVzaifSYcVfoM0Qq8M2c/XFDtWsObZCOnVZ2mBOxqwPrCLvL
Ao+Sf1dJwS++qyUAsnh0ZBHadxdR8Y8vssOXLbOijiDtaf26T4Z+GfLDhBvY9G3Ah0dNmyLcSBls
MSN9WeQtUE0itUpaZ67g/lT8VvY8DKapMxs+DYBeOvPeFvsTmetaBW7ddRfU2D4RiziEO1kdVUQe
RS+tbhfic4kI8l1SGL5mnt/SphSqWRkQfENQUkopGilyx131bvHdE776+En3C3sLcSPeBfN0yKxW
/ikL3mQj9iYsLv9QeedJjuSGJ4eAmDVcsPlpH4cLO/Pw1w8Ka5Ef5blyf5VhP+zC4EUCNeHdYxPT
NesRKbhyxu9zdZnszrY73xVgN0+IHTziRA/CihoUpJm5tUUubwLTbWCNN//yF8ff8mKz8E+LXuel
Dm00+nJkhBcirXblwsBAfjpQI+u8UFtY6yyyxpqM+RDTlwH1Ud/lTVB6LRlYK3V+/OJEm3SdqB5h
07vmrIzeJHmIIiu7vEq/TG8dXfc6tAcuVxf8yjDwvoNoE4YezKofp4hvw66GeljzAviSj2SPEIKl
e1aPTQT1BPl40lwUYg7ujC8so09/9FAoqhuS4sBwqG7lMIM/8DCRfM8puDdYoGldx3PbirbeKeZe
WREKwIgGmc9HxYkqIhIRsaj3OOa76sPsab4q1wtVnMkNdoNFRHBaJQbDDaQc2SDdxn20qneAPvfy
5X1MN9S0riBeAhJ8o5yJtNm65xcu/iHdtmUoNS2ZVhiiCBL0dQG2qymZdfRnqMnDXHgueC3sZufi
ib1pL/REweFm6tKbXJo45Znt0D4cjajGuhVO8GUlH+Lu6cnrGrGEwc6wT3u7penJK10RrE6IzeSf
EOjHfncouny6KVDtNkJJeDAJt+56sgmqYdv5ub/m+XplSKPOCVH8Nhz2wJu51QWV3satrSZjcjxX
Gxk8aE7tbI2qWz7MoBLCMgxGIMwtgK9JniPxP3sGkPvprwObk2OYW3l7HFO1pR3BsDDF/qGbRgmY
fWD6op1acQD57XUodqAZlD796y6cxBGmZ7gMIkAaVkSXtnTy4LqpzZmoOPAgBcp/XbpV05HaIv6U
DJGIYY2+Lr3AZqjb6CmECm8+mUMxJX+jA+dS8PIL7V09mGgEZa0nV0ESKwXqnlvpdbeGu+DXuHH1
iz8YOkfbD2tWlG9+Ro3c37auD3USKFmPz0ccozMBfv69sOKLKAW48/DoKXoW7xYEn+uKc64JaVaK
h8NLnhk8MPqv7+M4J+rY2tT6C8Og2Q+WQpG+XYvji/0JKOU0D3RlUEU4bK/C1R9auIoujA+RaSB4
B3lqSrDXmSPO2Hmr0uxFFWy0ksfzZtSy/jIJQ/hmw2nVHkTjRDJH4wjcG/27BJyEpUenNJdaVOQi
+gBR9ZNFoFq4J1u2sH3QyzxNPKzt7WtFdArZRwYWlXYEgnwEfQRxn5MHua4BtmbVLNvUcEtVj2gf
r8MRF5d4aHgJfFDRMuaETot2nc3AUPbqDP/gnHmYRSX0RdjIRdXbqMVsxXz7BbaK967VWlXKfdi3
AxRFNigfQhy/8QfvVrj6+NJjxp8ah/hr64oB142607hkJBIr/DGPYrnL+Z0i4mLuv0mKQF07upNn
RTlHY2xxRkVItU1qPpZOZ8VSID0Q82CFPDw1VQi49iCsEtmbj+5oDH0bSwKbcbw8+TMqw1Cqnn8I
Zoq7TJNGcjPyv531VMhi99Lb1y5PI+IeC0MLOtRat7RLxrqb6TNmzjg3O8kijRtZAvjS2GxqBJCh
jRDuekxU3iCshTEoLpS3cMV5Wo57Zk76MDLeqz4aaKhklNyTtWn7nzL37H2k0ZTBQF7aUizD5gFQ
yFOVOaKQy/6pF/i8zk97gSMtSLG5jTgHOcT2qILrQW5CyqrHk+wdw7iDPoOFv9kLfusAYuA4BlNQ
J5DYW4A3gbblj+xiOVYUnvoPjhwOtXb4F5QL2qtEmOFee6f8KRc1li3faETSRaEA6fLVo7Ftn3VP
zxFxUoQ4HOnXLXOAmFT14q5+e62BXCpti6ypHNtO8enS6r6wwwiypyPeLcGoxQy0VO3gUePITfc1
tGPGwGLhZAzPC82G3HMixLBZD3bLnj7U6S0AfeSmEQj3LzZ9P/OIFqFws12XambUHyRnh10SweG5
7j41yjhijis1NLAdZ4UKJUpxixb3CJJUt5Lgw/aYRKU9djam4jUDwkY2F+aEeoSsrSkEF/cochVz
0cy1CYF9D6boOf8DNZrB7Zfn57vQC3gQ8KUBcJyy5YumCEbwx1eHuXIaKfUaBwUbPQ2rWFftIHMQ
vmnMj+8dA5Km2P0AaupKYJYbh6MhWYgw81pUnlI75e9PHig8+yUx68e/qBf5rk8cBmwPWuQfA/mz
p4LZ3jptpvDACgK0VtmIM0pwH0FkXnxZjOvujjhMkHJ/hGiAVrk5wZq0ERTvYlfDeVZZXU5Iy3x6
oZYfPoQwoEPtRlX+TAR1l3vDMZAJfTe6Ie2cxYxpJV3YMCRk0g8SLxrC8DHbWJdwnxt/CmH8tAV/
tSMyFs+Ae6jd5nJZ4jdyFhxU992V5xb+hpLNyb+rnskUUeTKs9x022mDks0NZZaNlu6thNjzIMw8
OWS112iSOPWqzfwZ+skIT/ygvvt7xeCDsTULimG++5ETUuG2/cwKEohW1jwsfxnujLpUqRr5/psL
kC/lu9GhTeN+HaoebBiHdyZCVqynoaXdXBIQM1okINFl80L9EH1JMLqOY12xIkwR9rK2D6ZH4xEd
sv2Dt+yZ6/BgtJf/8w4WqlpY/PA5HrEeJOXaLtpqARrzNGuLrBFZdU9sbYxYYhtbZKyTNtCIU4/P
cQy8WKgMKBlcRH4Q9ItQjtsVyTXXR2PllsGmnHLusg0jpaoufOOmzH3mQEhSgWoiktVP9nw8QuDC
gTdv2OyURzHXXSULcfAmWGN1iu+Gw5YRXPr828CYDUTkXQPqEW4vvD1XA07uP3yztzuUvHuWbhTt
YbvHZJUSJbxkTGr7cISyV/4bKC4qfPp+dra9eqRXwhNYIAuH4dmfFgLysqR+icJjNxOED24EsPAP
jaQF/jB/gSJe9wzMa8kjLvIOtfqSxYLhLOWeYUdw3yB+62Wvn0yhgic1SMijlza13KxorKhsT3cd
DWq6qL2qcWwGHU8otBP0vGCnP5wNADQ5eCvEUA6UMXdrH5mYb4nuKlK4C7UASnYJQNX7xMockwOY
M9TuiD9PdfRrxX08DUTu15DTUAj/xucaR4QFDyUVUZdu0wwFlZLg1feLKp+ipZe0Rnds2uQ8SxoA
1r20w/8XWdqSr03yTR/I/7/gloasjySRcUb/dnsSIksi/Tj1m2ov1pIYudPUXsVd0YYSP0F9XSIU
3sEOXgX+r8WVpc0kO4QDRaqjCAYKRrGgGlKPH0KvvW3ENrVrLE43Z0pxAnd4oXKPe7p82SZ7ynGZ
Dz5RIjBaWEcGEYSJw17MEYXKVcTXtI+rvYzAGA98ISmLlcEV24uCvbFGQsTsC8NTCBZgi09cjD5l
KsN+YUwKKhTpBRhlAXAlEXyjaBmsFmh34XaDyIcNX73ay//wy4JDWJ0xeoLIX3jdYtSFChuJKc7F
T0/aXRQssHPKz3795mSEP9S4T1T5HQDoSaUkskvixrl+b06SKo+qNCtwbqdyBu45MlkR10QwUgAE
FHnVrfoVGXufTpKAPYH06EjOfxX4LRuIXXl1PHMAva47Yiu6lmktBIIXMgz4dhE9VjNG0rjZAV6p
pJ/B6gyu3kUnV/okSOShHn7GAuA8AudQuHsdueqgRqnsSTnZFupIl3Mp46/GZHvIpI64fOskeGr2
B0HQQndcXpcqvyII64OFg9xEUOIHPQznTFnZ2NQMnamsRGq/Bd6VAKV6pXoaJfnZqcG2MVSlWYoT
blDsuFLGaPbvl8XpniYMNa6UGcywFqQ5cCzN6yQYima4pURBVQsPo0GpF7buShqupQeLOCyTY3eQ
o7AMF8J0QSfz1uShOzoqCb6pa2L+XP4Ckb92W8yw98Jgorc8eCe4sdqw+6guGrJRdIXFQNA4/l0I
VKE/Un183qj0EkcIOrf7bpKZs7KAD8V8DT9KE+0Gpwop7JINQrRXnqN7vXBZPSyy8tocYEA5tydP
QSn3XvpI1uVdEQ5JblCQhCG9KElmqCdabUnR0wWvFMfdcOn9ydm2r0r+fHL31giBOUeruYcJ3F8c
wfd16isNZPpCyc4pTHjvLKHNP2DoDhYYmwvC6iC/fv+eMETTa47N/6e1WJ1YMWet2FUbHNpgZ01p
fKDZvG+E+LA/BaRaOeVmO4SYOTO32Cv9Apsq1ailgB90RAbdprL/JkLR8LuZNbE1Q3Tu4rcqyA2/
bV5P5rsHPal/XKtT49B7ukmBANdi0gTMzFQ5rf9OVEhe0jd/ySlpOLjNaHc+OcLWBTcT3B3xT0PF
sLgIT7HXJ7+OwvVeoTzm8B7LtOIEoQuQksqer9wWIwCxcW6EbxLIR8FqD6bRbQCZK1t9kJAL2vQp
MBP36eBQBJOEWkydX+rR1G2XkJ4EKlvGwgQnv3wgViz7aVeA8rKaMj38VBq7FKKdqM3lr4396Jou
YMZ1bwMqNys5exrAEolpfxTKrfoIXJuTvuNk3I0exdZTW6kdRlf6IhKouUP83P9/TpO9g24AkU4G
OnbmLuwNIf37ZP3IF6PmneOcPhgDNty3XdfD1QnheIL4x8+abf4FsCiOdM/9lAJrCgmENBPUOXfa
83vdbnIGIrIcwmttZZnJTmIYnuX/dG0RcLYIjKZ6/w8ma6LJQTUf/3WR4fZD3YugGxjhRtW+7+s9
WXP0WQtDHBB8ZAU3PLkpLD6qJxItN8rUzh0UlzXWvtZ8MvbKX5tRfMEbyVHAI4n6pKxCaMEhFfMt
xx/2rSdunqyUHHiOTzeNSKn01X/0AFNGuvvMRsHAEYhyorkFwTWy/utXCZPFRDOwGrY2PSw8iUvo
+3JfFviF92yLDPoQBupfHlh0hLX0Xw8WMzsbu3NPt4H9Cb0blbLaSmjlgHxm8Eax+it0OHm1WYes
YIRjoqdP0VRPDuzrbVx5PoHe89s4O68h1fez2NFwfVJfF65iCCSKusLvmFKbMMIZJDCLBOOGzxre
Ara9xI7AvZ4WQJqLWB27VbvSPiwZ3hs6o/L8zoH89efErAv80OEznnzdFsss7bQ55ndO5ltZ2fwZ
lf45KJXtFnjmkXifOU/lttuElzw0T3LQ4z6AM6RzlRUOcmlL2aNqUS3MHFMGb4kUFu7KqWYOPbZV
A81/NBev4lUAPL97Q75wHW1ZrmG5+SwMG9FL+j24KChnCLKVG1vdwvTrYPfzP4hBJwgnhK/URE8B
SFDrroqUaNt3WfFl6/VijNAlLchkEumB57xRBMJwBDVbu94H+GhgR2/w+MKE9epRROmHVsNWAMsd
x8zOsH/UvOyIO3wz7uAzEG9ZV6upB6ftl7R/HshhAt28XYM7o4feezk2bgR+mKkdkyIwzEv6O0CM
WUN7kFM/TcIDWSiGUMmPAUggBdYbAFuAcgDQLxxTVxVRpYFOPfxUiU0M9BlC241BgADj3qcJaoah
z7ocMZCZZyM6Bh4Ht7TZAnZPIQ5WaaWZqo5qq60p2OL2HqqrP08QFXTNdqIdJn58HGFWLVV5pbJ8
Ks1ewNvQGNp4VLaFBFeCI2v55MzdNLaplurhQNp/EpyBQmYN7kDD2M+dlG8KxGcOIu5E+Od7kdvA
Z+12DPxx8ATasXlq4SfJ0PIxKlkOEwW18735cphc8eTBP5Q7w2DlQOD/ujk5fhejM9thS8ckWK5J
0EwL7c1FaflsfSki5kmhpYArVKbsiBij3CwPHdoGBjR2SjgZF7VPLkuO0ArNTVYh5loqNTzwa5E8
Y4C4DoFYn8D54RRNmUluaun4F/aP47Is7imT4/hYYcDAB9AdfK0OBovY60J05mtnyNR+C34N7p/V
K0BPR2pvvHJsz+LZCkUTRn6FmR++mYdF+fN1fWveI9vw2xaFAT/UXKjXRoq0jb7ijQfQn5+zGXfC
eEAry27JgdM9RvrpFwwj2+xhh7cu1BLjGVXJ9rL4DQwo5we+UNpvP3z6JD6h+A/Em2lvzm8BP1KN
nVpyV9Wfh6++d9hmK3cpGTlMT99PGtQ8ycMxgDbO5y+gK7/IVOdXogKL3fxf3kKNRt0qujluX0L4
/pezTMxsTws5vU4f+LwPLzbZqqKbf7Ag98zp8F+pC370CiGWfci9Yqr8BAH+wZVccvovghVBSfhE
Mb0j4mN8LxZg8IwpyndAWiLx0BbBBv8WmHikk3WKbXYiDVDE476vNAETy7sJWeQRMKO4tgtfD02n
kbxCm3GbbMl1ghRz69XgQGEszMTQRs4voj3wMs2/VjeI78EIDD8VtNSnonrCGoKmYCGSI4X+438b
U5xgICWCicSJlQ6y+Kr2s79Ui1JHcx3Skvf+f8wcveZ9FuMJ/WwxsBIfrcg8zQkpBj5aoetfB4NV
vc0uCxPUwkl5TwhaqTSkwYCLhdqnAZUo93r3przRczvWa1AhzJqHjx1HQDdPeet3R1rfiQHtpc/a
6rzhZV5F9HEhNDV/zd04OQbF9gmjrfManAKPxRwEhxFzFBIUXx9C9sSTBRiq2Nwq4x3rPZBXcpPE
uyqLjABfrVDxpyrArsrN9jfXXVu9tOdkM/G6midOsjTpdUz2E8A3aUZFwesRsEAyRxB2xRIdo9Wb
Pru2S/V3V8FHz5bhhS17S30TJvYj/3IZ51qxQj2PIGYZo32zgFa1cbON/0mURKJusBcsPHYntRJh
tAb2vQCAUNB/AqocGDawIlnBJ+gGP52B+b+wm+51j15K86Farb2pxDT7HYFglHY1u15QT29qM0xp
oU1bL5v6tThVQvFdgr47TYdIDuMlsu6dwAYeEkntwlkqRP1Ai4Kne2Wrkyk3nqdUxoEyGw9XC9+y
ySanWxFuQ3F+M6e8AgRTqhOn4/Lyn4x0tiHlzXF/M/sNgMnyEULvweZhn88F1AzXxES0C9RF8zWv
iXcE5bD2oKjXMA1N9LUW+W/Y3cke9aAt+QQPGfqeyh5hh8HHKajtyizkXyGixfFaDOVL5T5jo7jz
QGQnzh/BGcg7A0+yJgwnraiDiDA1o34mHVHbstiBLaLlOB0+U01mHf7SOU6iQ/M/MFNyNE/ejqwk
ieaDNiXpSJBkHBSYVZEM+ajz4pWQQ4KaU+YdtUyifzaPGEsoEa6fKcbeuPVW55RuGwChgqUKYuFD
JS2o/we5gqYMvoFszK/yr/QWmZO83b4kzlzBV5vN0Yk5KSlH3yqGq2smhDK0HyLqdwJc5saXIPhw
C1h0KLMSu763QUK4c0nVkuyuNVOPWBH0ZKW0/iEd+UcOSY76RP7ddar3iIATKEGJfvBMjywSLA82
q64wouGmQKreJVG9E83HK9UlT69tw4MwA5fuoE5vTgP8VTyvF4D8PfMupmxZGSd72xfE786XvpFX
BhkZecG7eCXqzYN366YDyR6qKFD1jPQ6z7pWalAxdAMVkTYetNED9YliTeiexd/VjvBg1qpG2NGR
NsDVYGOw7yx96iJnnBSMHLfwN0Ms/fxSQyR9do/3VzLh4DJKUCAsqnmg+i2r/IbG4kJps2045F4v
Zq661V/OKifvy2xNUp1eAK933cV1hwdog3yVCrL7bL0Jct/DFZO4dxzs+lnSLOX74tzcrLqkN76o
tdqv+NVuYaofge5QX8vFi+OAA2/NNxmh+I3PZXQbrrGeKwH9ETFaYn6IbIwT+XgnhJbAmAJ3n/TR
CuChErStX24zZrzZ77exfzGwPXZ7/3JLR1/QY6Uvu8B2FpY5P5Kl45uW0iOJyz9DyHTCCkaiLxLb
6lKA8KVRAtgkk1JphYuMtEC13papYmEVWNEHbPJ7kTQAnyL1E/CscGpEn4rnKwzxim9Mqg8Q0VT3
S1oM0jIv6si87kRXsOgxFZUG+kPIDJffJT81HKDYF5621tPcHvsl/HtZk5TkPcTwVY0+Qu5XFckL
kwk2Gp9c+vikD4cW8YPs50j3ISU9Lp7R2kiBMpSXZ356ocd/pTGcBJDsUpwsZM8wk0ZsG9gazDAV
C5VBIpWlq7EIG787/qVoh7Cpvu1d54hre6vAzLKMByvei7US5tFQBU/oGdnuxcK4s9jYNz3dyUGO
43E9l3tNKMBvqDFTmHsjJf/Wj2g1uecs9xUVbtD+Yoe0+Cu4tV8SxBnKLk9kKeoEq1KAMvot78Mj
1tdZriOj6lknZ2WtkR2wtvvPVo1KZMwv4+ZcoqDs1NiP2sn8Elhs3w6t6533KqW9GxQPboUoVsCR
u1+m+1WGzASMPzTcpi6l/4Zu2splF+qYWxRku1ooE2i/1nrO0OmkAc1cJZYp1Oss4A7kAz90PCCT
EvvRrcTk/3IZpU3+d2UELpnwPOdx/hv1cw4Q2i/uO0AnPfwvfOTtMISroSNOORkGnuTIovxSKsAk
Q6l7KqdyIfqWcqqivHHTnXIslZRZ7584NUO5hvfi6kWtfg5UPMZY7EdOnpm/M0VaACiXA0lPuWFK
2ooxRTmJh/vxlfOaEa3vPEJKImHhe9+EcLnp8wpmTPseUokAKgd7Cqe2L0nMJbgLJqQHrAnhK+Kv
jeyikSLgGUcrl2bTh4rZ94dI2wm8mWVCZ4hwRqqiKftsGolPDdQg+V/8V5OTb/olwRAA9/4kZKe0
8uT6gZXjxD6NyA+0btepfFBM/Gzsn/1HoVDMHNp+E3PxPX+7e5tmbQKYb0rEpPWkWGvBebUx/dI5
0Psqvwp1HNLk0kSmbj1BFJJIVNAozRsdixCdKbycq93CDSG1XWkAWG3y55A1mdab144LSXs2czd5
T36ceBh6TYkCuToAc5kG6JABwLlGsSdxsa2mULy0bEF4PHrCrJDY5xMlNkwJ3mgatKmuDgwZnehN
wKI9fod1gTdDk7tH+vkessxhFq7Yl7zUIaiWkdsKTX4qItFmvWFTVsnnuqCVWaC0HDeKDHxYm16V
l1I3z7JHsj2DHSf1l2y5Kvac14OXLc0u4ebETXxDwGdxOO8ejlOTVpN1fSWsnb+w8ehVsFZD3Ml4
XUKtQJ9gdDHK0/EknsjJOoAJv1QS6Iw3SZA9Tp2VMuZIzon7krhF1eQ+OqLMJlAPBnMNPRZ2Yq7K
w0F/vHVqIVP9s9F/u8bABOcZtLf0hrl7goynKTHzjlQuR06RdvQ+f/zT4v3zmvX7AF13Okw4+h5i
NzaMQ8QdRmLPbfZl4WHzjTqhYS45Dry5Wfw4RZapqEs6l/VjSkdXvH5uxuopPtNwx/VOTXaWyxm9
g2JKNiCEw9sfnmsSYtDGQwJF44sBMkAXoPaaMRw56EXrZO9QmKftX0jX45uVqCKfqYFia/PRALb/
wz5BDw9lxOaJztXJAuDEUVJwARBvob5FgPva8thfLuc1cRm2WQ4hjURvftsxBTpuUhh8aMURl39J
7olzQF1vQFQR4K56AfC54q9e3+tygXuGvPpj2Nq6xp0g8iyQFTTXrvxVEiVHlS4o+aubSyxfVtcO
IQGPUg6YJUm1J8GdioWQN2d6uh88A/EMwTL7FKTQEeSLPuhN1llscvwDepmKLzS7tBEeRa3M4Dfh
PWsnu+yIrI1npshgkJ+Ph6xuVe+YC60Qzu/4t+C4UbDUovhWefrej5zFjeldG8vISuFUhhOdWzo8
iq9nBtjBPC81hlXTLSEUhSH/nIY+mTjvK6so8G+i77nsQ1oiRR1kEHs7iAJ2BX37GSBmhY0e3YFQ
lnj9v7UdmA6Uo9avSx12ri0QadKXlFBSR7HUIdYjW1bd48LBRAy9emko6XRS+WovtbSyBmcQTrGq
14aS9LQok4WEr6/0jlfxgaHQlN6/hV1canWpJekA4fzvfFu198jO2PyMJs20h6K88TimtdGFl2Yg
ujLo1ZgKSQplm4lfsNNdDHsd4OV0v2iioeAD7H+Zo23pQXuEMTRDQw6gXnlRlEpqAz7crRXBvfYV
YASrJPFlDuqqrnpwiGRRnbGre12HB4eYfNE2vNN3INSr0wIFQTDNm69ChDMmjqhJEAWijfjm7dHk
S7NUbaHLWUhzH323cFYEfKRPFQhLfNtKG7f3xDtX6N14jifd6O0MoBa3TzZxCxPhu87EXG+VQGOW
DL7DRpLXjWHfZf4UpxxhfgVUVp/aAFYrrfglYj2OXYYgnNCNXoFqpSbl4TEg5nG9krprW72UBMoH
nGe0QOBcXXErVdXxBtw2L2ee1PMVv8VKrLhz9v/iq4zByVEaRCueXWllwZAsNRq6ezcPhoyPcEjj
E1cBWaoeOMQEj2w2lYC9ec/LyFxpKDAQ/u1Y1etgLgYpYnW1n3NTvY4NhZPBZ1c7ZGtmbBTorGs4
RLi7hkZ/fOxutAx+bMhYvRnnEb255x7FjZEuv8sQsVtVRTIk/ACDKLnSTQ5JfEUBfCh38WHMQjO2
M66Lq52HjtUd74Zey9B6O5jSaeFUrb7q6p15DsJwqlWnoHjfU9WPf+xF7tAdkoU8KF2mcPNyWQf3
M9yI2LJ5XE/r/xeaviBFQ8doIMDWkAjJbzv3TVUCCneYDaf0ophN1X3APr6owYHCkNkdM8LISiqp
Y6Imt2zTxY1+86ZqScBD8lUk6rzjqO0vS6GhvFtEDfWNZBhpKc+2O0bHv9qXEettYy82uTDCHUEA
ArZmXmt3iBzyakFBJmA7yblD4yJRrBhmGsKYc680bzE0Ui/LVXj2SxTvhHOaOrTuOF+v6UCaqC1D
1yUxFRyzrZE9Yp7Tiw+Xy3UARO++GDOX0RbMhh47eWAbhqRdCCFXl2pjN8eh7Gyu/MaVqyPS8BHM
C/tfqV9qs2mYvWhoOrWOcn059ayERVbPEA7+/QWctFfpMZvYuo1zh1be8yJUHqHhC6b8ksz6+kQS
Gap/KsTJPnwC3cmnnRFx/QooD4FVGy6v7SiTnAOSwVefqGpSFMn6+99xuElzSCdUl9Fszzp6RhA1
8aynQSP2Jb+3XPzb0Hp0e6/1XZD+iOD2bxYYNLP95h31mEooZ8irLXrRrGkBrc6//1ZfMUkP/Hiy
WRJ7Ri6nUDOYP38TBhm5M0UpjiawTkIrLJOUziefSms1yECl7Va6EakYoFsC/TIB2gMHRw0BvSgu
O3gOuymYNkk2EZ1zeWGGcEVeKGNM6hDA0nH6uldOSA0dRJ/N6ARX6oF+n2TZdcHonI7tVCbqkddx
KoJnaP2UvEbtOMW8T5RgY0NrSd7ZlExTqWeYi5dOsSED7XXBn7JiUMwSxCZ0te/BJcaS99BpV+Lt
vIu3qpwhOaGhTL/YIhd0GzGww/syIm0YIbvSk5piypYEXKIQiVciHQvUCEAi/WaQ7wM0khWCSyR7
1HwT/XHRJdsK1jAEyLOuDmLhLRslR4sbMzyZkpH7rw6AiW+plTXIV4w6+aqN+Wel3u3ZlFlGlAFu
XGJzxT3VNQ1wFhe08cgtLF/lJ4Gzv5ruCeejk4N3mX/In7ubihMPhAZSTmE4Nl5Yw3Z2BpRW9MWa
/4sB6bIUNby4KJ04vCftXsc+X/56a7e2HLo4qx2gLmnpUUI49lGwxPhrITZhUd73AemAR2Xdbw1F
srSqEvI+1eyI0EzjmFSYwUKKnklF4i16hQObQRpaL4N4bXoio3cU/VUJK9sAHARIgH/Z6DfXaz7r
MA9sRwVQ7CMDswDjwkLpoZ17TuT6Jn9hc3SqfwOA8HbUtdxHuOLmJUuz/VeoiU8aDDoRHUBD9xua
qlcXRdjjBFxx3gVJNHiiGJNkiXw7upybyCr4SoUuAk6BfgTvhhwaRMT56qSK6P1o44E076uSHbj+
gpR9VHfrzEnVfGKK/7Ejmga8csFZ6V31P4qnWh7Ni4Y7X6wb4YNHyd9F4pWq/bTpv/EGdF0u6XUB
8EjMOKbC3/A5YAUN57nHTTqTQ5V6tSbVddfPmPrU4op9o/DpcMklqD3lxuzvhooKT0AwllJXe5hp
NtYZTPC87ClaqTURS7XacudU5eor0se8zJnTKnz7523Cyj2wJLbBv1a2pss0pmco5MFIoyWj2z7g
/N/JVCxnZEm3LEU1DkwW7svaQ54h2HJ+pgdB0DWq3MLxBiMYNonClf81lybzXI5M3DihP/OhO+/4
yT77aDK0yAaduOf9e9ND17gdDmRw+9+FXjN8j2fTDDdLly3eE2psfOCoOboT10Qtjr7RM9TAQy/P
hrqkKrClVJl3g9nXT0wzk9qYAuUW/BP9AeruT///TamDsEOovLXcZhIkQ2Yi3uc5h/hPOxD25JMn
edTxWuoFykmMkA1pAPI9EplpS4QngPXKoF15NfLM6eJ7SFING/rY0Lt7Wh4X4PP0MeQWo2o5zXNZ
q93bE/GPJWWdqWaKt8pn3d4mtTd8HKlWORrCbl4WN4IuUO32f79NaLdOvLATFUxQ6TNRnRxUi832
TIGK2X5ix4rAjZm/3U9Wnje3CA8MTr1pHQgvIAQZkseuVQWe7Z4IWXVuvavhBn9whcQzHCm76R4K
D89hnLsjGn+g4NO12hnvvXOrKSqVyV97S7CK9Qd1OKEfvcE5KTSEdZUfyDEd3Ar/McDxsh1iu9HN
Q9mDTS2/yPmxWEqwfSd36oyrO8tKr1dG8N6W5Jye3n6HONsnpUJYtiwqO5fKzYDZTxgyB7D/Qh7b
zwnJyd/u24r4Ns2eDwkwm0BcojveX9SRf4K7pselehHZlolg/BEFslPJsPjjpi3MFoMOKv2QTz31
DqWqvmeglfmfOFfWt8TA4jRIe8Zb6n9rcWZd71h+KasuFQJbWSR1S0gycFstCzXUSWNu+3d+Kujf
MAs/Fh+3zAIDoZ9ZRGefkNLPOzRjd8XY5/xvPAtkTP6CEsgemxy2Q54r6DfMITnc0uWfBq9r5zEm
gwz3X1/MPNmiWAqPqZ2xSiRRP1UG0UGujF5TMhA7wYPgXDcfBL6utTPIoybbxHwpT7FcJyv1X6uF
8ywMuVyfNTembSZcS2aNuzna/M3wgCGtd1YuAU0Dzem0rj1Y7kdFlaFhNbIdulnnC5TIs7pdohKq
TS0AjTAV4QQgpVr5w/RdEoILk7xFhoa5DqDjSkqEAoc+w4E/9BMdbMDgaopY2xiSNvvz61XkcH/n
JUh9idExjLnwdpFdj1K9bTqHF0gm/ghjH4HFIF1F+FpTHz0utNOQEk4iOuIvN8xOGAGZKIJamxOX
0iakmrSrnnPJBkCwRfT2Wq9mHfyHgirvlEXR8qL8vAsZnt2+DQnFr+tH0PLKTsK5yv+y3mSt6JSn
gW9tUyl+OvUVnmg36HUZPJr/U7p30Nok6cscwAQw57VjZkoDtsA7nddOhg5q+IGSxYTHVFW+RxE7
BGoayjaD5M2so+6aCzGEa2py/8jDnDxnWhPi9d5MOUPMCxHlEoxhmgHUeQXliprpwbke3meYurtQ
bIRq60Nf4Kkls3x84AclUuvCINFdEHWCtKjFrAQRUCD4AgOchJ+/1amUMNnrSyYc95GIeFgxDW28
4c/cnDuYJDUMKTN5Xim4eEClUioFjTktdMP64BqJrWc9h1zWcrl5i0wG7bq04JZHvfuiiNkXABYK
lxlobGfwuV2jKNlgBHMb8xUv8f2hkEuwqelRIShzbOS9NlpLKg7AyAXAfIsJXlpT+DW8NakRATfb
hDbCKSpCSOJt3lBye6hrL7twun3WsyHihUGTClAlVrsRzdnwe8uMjXOf8Zj6BK7umHSlr1GzAi3R
t6UubOvI6lzkIjwp2P3IPybt7umcFjsxwdADdpuDkrhgL5jkRHHTlkKgJVRcScih82EisqJI5rrG
24OokZwUih445G6LuQEYHZjXgDjnZw9pvGlM+XM7HzzSvhqLPfWAdz6Vu4WNCUDqAlyUQAsoEGRP
3CSaSwQ096scTKzZlHX0n0V8jeQWHeiXo+6qHFibq7DjC8DswZRRanYbf5g+AB2mcGUcfA2Y8SBV
cyd1webCNNnB34IOeU8NyBzOXY5On6LBjJJTF46x40XrqsMULm61H74Eg5l7Vt9d4NdNJP2EZTOP
lKXeMHti6lhDdiIFlM3tWRXRBdV3UeAk4tThxlzNROYpv1nbSkiRGk3dWhuSLIHwnw1JUN9R8CYy
Qc6HTppZsgLj1hPk6Nwb83bzD6VzCi49rYjMV/6IfRL/yODBU04EAA+MLU2UfJ5ts+ljVMhimd4t
qZ+COFwAnzyaBrBj8eF7OtA4NqQrD7XpucmpmhECsgnUHbIu9VidqXfcWKT1jcA53ON2xEf4nxvO
EUtIH1IBAexTfBXL1UFIcOPGxz9byLTG8i9UFG1OlDTwwzzZn0CDTnkLSfTL6QNTCAQfh4/GknnR
WUyBaVJUoQo/k7fPmZMWDPopyiHc6L70KhHyGKnxlcnXQJ4uJPIv8ft76CakffLeJiSDJAiZS5CN
soEhFcjp4j6q/phuJnX6/p3UbakEh31ksfJJPaXxYNhSNoIijcef+DSmzJa+UUe6ilJHormnBw64
JsA16iHFIs5AHKxDRsH4spirP/7OHX8gXQN8IqPKzQPr0B4S1AptzNB/MjSPGGfpq7pqMCkfDe2J
Patojvgvt8L2lfn2Zu1sL5zF4Gp/w7s0OaUjOzEMyskyZybPYq86MMxWRHqIPNUDJDogeeLb3V2+
aatu1XhKltFvTdJo4Taf7M0Lyq7EPiRb+72Rcs1riXskuNTWx2qz8hqYs+Y8vYVSsLy7hOurcYAD
pWxyXAAyQgGpNCKywLiX/HX40pVT7st5iuxU3l4De8dp88s1OfiIitnZTUrih7R0hjXCZSm1XHqy
D/VNzVAZwMPV6QvXF9uIenF4quNNeleD4RfRbseDZaK97SC5gh3hqsFpfbHj96AUUzL5JuDbNGVw
qEpoEA8a8bPR9oxJJ0qub28WB+n/8VCiQR5sSzC89UDv+AbKGod8PttgzbCIrcX6gzADhjEBEmKi
8okEQ6U8iTLjnsOmwUmS+lWsKebjNjV7uDxfOfdgBip3RVU4/w+c2akjtF57KlN7yZ25GLeB8sca
Lw3o9o8S0MydNVuU58c3VZrzkMz9pJRuAAOTtgZ2680E3kKfrqq65MM7rgLhCrUkcAGcOFriqGJQ
gpknMA4QtVi8E+dO7BuyuwUpvXqr1ppSuFg/JBySJF1vERHiZOnJfEE9vnbbnIL0ms/LjQcIsubu
sa0l4vjDTRMriDdDTwV3pLA+Yjk2XmueyRGwAbnY/U6zDQCiKjhMcHbNSlqJ4b43WhEOTABRqAep
ew6pAOmi+C4ehNsJ7yDgdbMBOs0uFzmM5NxJao4Q5lofRuZbkZakDPPc9iqyf0pIzWpAH2DTM4+c
zIW1AgvnWVD6+J5SP0dRT9Xt6sJNqkgIwzax/BZMN/phB/oJC2rvCrzi48cprBxj8UhYoW7fy4Oq
2Dnl/xzIocf6OYwczgGlFmEsFxIfOCCmKDh5e8aJRokc2P+OIxEiyY/cSxtcdUGj2UTm6D6sLibX
/sRYnlcZygcvQgx8eiouOlWsZkWubDq9au0n/YMI480qFW1bZPBlJ6Y9uL4OjrJDPIwWsRO/uAlW
g0KpeZp4I2e0t68pa4BThZ1L2QqjLNdveSa8zg5ITn+HA2/Gs2II4/3QEagIiDDs8q/gw2jRJBA9
b8nDzNjMZpjRKs+a5oiqzfRHhVbkfQoXOapsc0x1ICfbrJ10zY+1MSkyxDOlR2OqFzY9FcnRfPOg
84lQ+zFOBNbcP0ZUjKAHd3cCF3g5NzDkK41wgpdKXYFNKEL5oirM77qkeI3UyRdkbk4i4CDv44zw
chaP2siyz6/rIxKXq8Ir9BvrM/Wqg7xk4JEMe/W7f8/VP3Rox9e1jhbpwT4Ydb1Wdc6lxIGs93Hv
kZV2nTT2NL7K4v/usDdhCjhxeJjYcyRMVFseQtEmb4g+HuTl6qCOS5l8+Js9lsLT0iORtgdE2c/b
uRvo+BzOYpcN+X1BkNr45qKbW7coARSYPBO9BLHOq9PkNq1P18tu9b+9iTfs99/U+N6AXj7T8E3H
2r0gAVYR625f66Wnyg628Jt41Ed29/c8ZNjVnhOiar9IqcEi/fUlY0VaMYgZj7Cz8m+rA9h2HIQ4
c0SIVvJaUem62uppOyAXz3EtkslcW/moPkEFXxnB+sNpOAnXXac0KpAA7pFcMPIQc1t+Tdv/lGqY
cYbR7xNtVquRyGqGZBwqBtB4MkzCU3TycHfzUCHD8bVAHYMVayK3FLHiwcu0fhch9nrS+LevJQhk
BGAKVfbd9Ajd8jxlyLuo2re8ir3VTsGpZVvNFTBVUEj44zZ6k1I4263WNeJzOGtNrCYKIQbX47zs
pdjqOlqSc9kfCdDztKJVGQQrlEyCOku9PqMVoZsEFafPS1VMjc1osAQ9gB6beS77rU7Q++OXmfVZ
BDdVQepMTm3AKYGHcWNnKWp2Cz/tLdsOeNSWZMC1yCl+YyzNW4vfYLaqP/Mlrx4bWX4QQI9n3CjI
sT9uLTGFCCvKlz4+1rXhGBb8Y1V4GfNhrHFLe5oKMKuou+lUaFlpnrE7x2TqGn4mg1ESk0TBjgQK
CA07SnYjF3o/NibjE+2WMltYPax7BS2GrqE1j5bsEHGsxILfyAuLNhRgpzzb+XM5bAyq426hbBpv
C2YfXRntE77c8Hi9iHLZ3HHoCZx4K0/AMUd59dSf/XaRpoRnbzViMrqYy0GxzAvNlMQ5fEBVuLvk
MUeS0e9PcA9yNi/fBgyUKyMLjOPXom4HRC0vuebyuB3rvzcnInITUA2XbHhrqN08bQDreLhirBL8
/In4MgTutXOfS1TawdBc6j1nE09QvXO6TIPmV9ZCdlqXtvB78p4SwhR/BilLoblsJCSwNZEL/drX
mHIhyh0SJqnYW0iXmTcmN+2nQQvDTiiF+N6ue9fFs+8AIHkh6BDm7JTBPxvJ65W9VKDoqrfvpFK7
j4E9d5ocpY1ZbsgWI774oUUpPePbuZ/mH5S9eP2ugC+xbtgCrDp2CX1/RbfRB61leN5dErrKJvkD
a6CJv+vndJF6WHaPrjLbnPSLHYKKE4/cpLhcQYvbDiDCp00+XIg11fS7Lx2DCAAYh0eBTa0+7cCx
oVSqIygMY0L6d/qxpqcF6FUSxroDtPF+C/IQ8Q7lVN0eX+ik1q08sK1CxfVBXNXdPwZb7UTmZBOZ
rYMmBB/vbLuREAmhqtTnSU7EHb4vojfulcinqVPrOSCJwJqDbW+Udi0I1P7FxRNaFodAqfN6bVWB
FR3/oV8P9ObjSqTnifhun5hUcveYdRRNq7jfgmDQF5SdN/i7NwCx5bcKShEWDXALWnclEUCLqIRT
UFb6OBVyT6h89rFYD6sHpsa/FO4Ss8E8/2VZ51XGQf5mJLS2ELm9TvgpoNefeRwvD4TZyuCSaUiF
yOlVGcVATJ+HzWgnzrSpc884EssDX11/CHm2jZpZHvDSEnxqmufQkAtg5N2219szcoWS9V+jtR6e
YW0onfIqKE+Vz2kiSD29e8Wwd9isd05ILX24Maf5NiS5NnTakXws1Z/ry9dahMT6zSOESiJMAIiV
6ah31nJnis3HMZRKpgDGC3eQXLiGRI5TdDlzUHPgWw75I0YnN1k1FdKhWXOw7nsZ4XFr+xydsptF
2lI8zQ85ciOZoHf59FxiHSNBKw3wf4aKsutspocL9eH6rEHt+rMkBa82zOBTPR+qTbOvBMOYsVrs
U+cXKuUrNrVXfqxZ/7o3l/TeA17+24SCNx5DKaFPxGCJEUpTDC7NEuWz8m0St+o6+3XOrIfRBjwv
VnmNNaJu/VPEOmGOJOrKBFEFYbe3BYScGXoWfBrZbgQhOySMG3v0e4MPMHq54Fh/TnprXKw+cygV
c4tYTly4QTdvZ9rcb9AlwuZIlRE7fNUXhe/DKYolB0u77QaqPKNY8zTUxSA0+XlNeRwxkQKX7eUY
UVq5ngejFFaxZbzBC4Q1s6W9VRClDvwsgUigNvvDoIUkcFSrtMHk2Lgv0HxdzJRNRO5gJnlmMr84
osektxYDoJQhCagslSLVVlkn7VtSsaD2qWTDsbBIri3/Kd3Z/ldVsM6hiWGvoM1BeTJIdEbfZFJY
1T3DS3pkRJTCCjZ76TXzFuDoXPOhyeDFG04z5jcrbdL8IpQMUg8Ty70+uyVHIgrTpx8Xvx2z7DkW
OC5LMStQN1/IYKgy5qbB0F3+WuKGncZRiAyTH+8fbThlwn9V0jxX4wedhVqy4Q/TDYacr+/GT0i+
/uxCjJVA7mu5tfoEPl3gsC4IN4TNus+dGQNJWleFonv8oe/khDOtbe8Gth4or1dRKpNwz0LgtdGn
6JgOVoMTlvB2l/N/xspuy7eq1MVm9YtZmER5fNlDHutgdsy08nR9tQPrSQ9Wf0SlgFQvax9ejbWB
sEUM9FXTYJZVnIO8D9fw9wis2E9SfffzBsrRu6CCPNAUlXLh5lAUt88piC/cAETchu6duPP428+4
pSAp6u3TW8ZUGP+gL94Wi9cYys3NTEyVqQ2r3rYma7/xpkWhMIFKxsOXcDxbeVMdNEyeUFmp15Ix
xiqPnhyMGP88C8w/HRlBYJ7D7NguoSvW/97uum9D4Fmd60I5Q3X/n2jVeX2USGN/PTDZDIIPMgz+
Sn2oRLQC7ygbiWjQV+56cUoPt1JQEwDKwBa+3wrxPgj3SMafP3u4wib4/BubFJS0mrztcA13plM/
jVSOzgooo21CdxW5fLeFlMHTwDWQo+DYuKcQ2IY4GCY7ZN3rc3ksQBuMiteYXo/l+nG9NNOAuH1U
giQNbD24fG7s5oNuZM0CbScg9z23JPEeO1LE470/eoq6p8GHyBhXcczRXGWpWtzH/GFImASn9Pcn
Hv2B5L1ulvHvPhgu7p6hRSIMnY6zg5MbOUxpvW+9QWdIh4hEDT4aCi0vyaOL+5UHUBu2hBixG/2r
/BhPnE2flwsBvncQWXvCFA3NvqMjmQ44xfEHnfzeb5K38SsYtTI9HWvshEM8tjto65GSz0LaBZBF
T6i28wkRRGoZnK57AihOclWdFn5/ZICYGFEl/RLhuv4wOkLhyGWFwuIvfCl94GG/Anj+tRZvPHEs
UiYC7MCPYEZqgRPnrN2ReBHedos5wf6qQsYfF8aqkvCavZphO3t/THql7UCY63XimejJSCxvpxMU
VXvuCNPDvxrTp3gwHR2Xz/XfX2kmpcb/d6Pii1pqdBMIfOizZVvNkvMjU/Q+GKyeNV5Q/Dq1sIXv
UiceqaY+WxeWGrEwMOrPFvnFtxMOelb+zqnDlIVRtKYkuRwlOa7qdi74NXy3YOBCOuE3lLoFLpBW
oPMQSww3dbCBxbE/C+cZbNr2JLZmxSQczt2ieXxs5JQ27Usv3T6hNufLqBlkyGq4qSSMSkFzIP1Q
6AlzqGzOgr8biRR6PMc86SnYefIesbC2mxbEslRHB/MWcyCkyymIxY9p63vCi2GfrSgPdkmvcyjT
B4LF5GCAf8s7WuSo/+M0j2gFWZSiR0F7czUf+ZV7hS7b4oWINfkVDIAGnSaihMoRAVYaPBwXiJuK
FfIzftObQ7I3VqyvhuHXnzYTRPXack3BlX8LfR0ZWLh5MhwZpcw42moOaoIU61PfrYAPL4BcSaNx
xuq8LJGFwB/b+vRtnQSmtoAPAczhYSFWGYvPlo2Bu1zLG6RR1la11xQ9A7Lr760rg1785dRiFtX0
2ePKVcMsD9tA+iollU1Nytio1ejDZ+QHnR7V4blV0LBLPk/HULuBL0DEzoK6OlnxCxwKhrGTqxMW
SooU2bmYdrANSu/R9jQB2S3nbOCU8fI9uZGf8TJs9Aixc3dE0MzshEDb+APYlp6rp4tDjqHEeGLz
VnqEMQQyM79ti6yROKjC5aLzunJd6cUtCgxV2Iyhqa9H18Tkm0yhA/iOgKT6wL1TTqwI01WmvQBu
M5wkbtkAcSMMUCmDR+2UbIYh2MurMP+q/od7Lns451RpPRUg0dGQ0zAqiouXiWfXYNL9YT/RdTXB
2qzQ8tsgDn+hAmX3S+IJ6MUxkOTXzHDBA/Rv2ficWQNJWgCiwmd/W0hulMD0hVXtGSlnpfJJ4rDk
YvcP4D+8erJ4i7mE0GWot0RS/1cbBLMBWMZlIqlefeK6NFnvqwq6T80dKqkvIWo56udzbwmHqTqE
JWfzjlvzu91VlicGvIFrtwTNRS1jA4+m7njfRHBPc9nQ2sZ51uXfqIACV/KQVdBrXXB7Gp8P1T5P
S/XMm4h5Yc6A6Rdt5WRTOkEWmA2M9KvHos1sSYKjaiGr1AzDwjPgWqlGBMEd+oqpbg+Y1wo3fq1c
9OLqRwKqiCWjKVnIKIwI7XWVvkLRO6xhmKaC/fZnZBJomzVDxnEcVqVY6D4T4YVAENlVJSxC8GWI
86u4OGl66BMwoZ6Vig7ASsG7Qf7unfwjf9cUzQ8tODaU/RhaZE2pz6ttQGWNvYyYdb5i2kiWZ7jl
zLSbgKk2BTZP/T2A2rwCAmiVH1/hirGTNIGV4nF6mZTWpTrFgi7QlJpquUSwiq/0f+jG9E5r4L89
9+Q6dLP6+STOH0QRi/nhVLqu3K1RYwYVV+xVtqsZF4EcQwWGVQxdKnwWibMns65kfeZNsVLI8vUi
2gtvkcsc0rF31mcrnlYo7utOgzuQ3wd0mALHWL0MyEEzWomchi8YW/pcTZMrNdNt/w1aFGIRcQu9
Lj6S4YxmO/z0DcyfffBsypM6RizM02b/VvMni5pPb9+UNN4A6h6bEDJnEO31h3hhr+dwX22HqEnD
pPuJ/0oB+3Sc8eR5WZgJ3J/Psk0hwegieIGJVBMNnHbJ9Eo90w3OoAVRTHXCHLwvMj5aJsWGfM64
nrTsoL+pNUDUgIrD+bWGUH0dP0Pb4rs87afHlcbx/K+lm+fnsux8k7NrTzpdWPfg/5LnNWXgng5n
ycf/T5iCTvSj1xKS1qVL/2LDQ6NO1Ng4vizE18e3v/MvHigNTLqjmsLbK2PyMn3AXEGKOG/YtI0L
V96gkA12lQvWLjV9VcqKGFiaKgi1tnBifNxiB4V1MlPS5tIn1JTtSnTUoAfqva61JzFID7r+GmNv
apMVaZhC1ydbMNP66/oZfQ29EJFjJLUciA9SHlBR3J9lWRm3W3WXees3+rjLTh3y0Zg0bH3yU6w4
rU7CgSxOxqOplgvJROy0YQb20PeQHFU3Rq6ihhmiru2rtf2rWdpqJOf0tzII8R62NvZMAh+ywAo2
pRVKncxyv0KXnOJAswH0zDThqXKXoabTV+QDgI27CX9nEjh8EA9FnOSR+wEvEZ/L/Kh/0fkqwZLF
RxlPUGML4R9ntLlmSHe8GWOVC/FiAgDn796GKo1CZs0dlNO9XON/1E4I5PsTwshfYQnkTFJ01tzr
ofi2WHmU4TGIKNphaoCZuXXR8tluXbybI2GMKEgVPNSqiQYCROW0cNm6dlL608n5CA3f9H08Dofi
7wjwqMzelegc9tvUAB4+AVIZJKyy6piaXySKiAzZTQYXKXRQhLdIaxADhfg8i6LoH5p/qzfaXTFX
NtMyw0jJJRpnC3Y2uXMYF4fgKEPVPZvW29jcnh1JCOfhkD5baSo3ERp9R7OrpQnbbUGBW0a/ZtGT
JObl6+LuYgfdDX9dqhCyDdQf/8lyIeSHaGgBi6Xg3arboapg4fEUnYBQzzVqGc4iI70KwrqGjD2x
PHStMwuC+oZ1hToHkstBBmJiVAyAsbIG/U5rPLrEGPRCAQxwu/lxexwu0yKAJbIKKW3Wiz9IKBFU
T9obahbISZLC2vFdPJEzw1saXSe8S5zkaNLDVmDR63OvXz8CU3/CQ/WDictkBdraAoXgskMbp5hR
UnAZB+gewBkJ+vkwdL/1OJasevTurEok6txlCjI9jMSt9Dpvz+ELubu26el0Qp10oug/q24Abyk/
FDvy9MascTHajvf5E7Jxhb8J+pAhEPAhTk/LhF9zckPaBMNUf81NUuF6QWpuRU4Q6rz/P7xgpYlf
+GQ9G8Cw1o/qgeEDdDbvs80vEf75CvFa3p7WkdmzjZdSVTXn5Pj2ZkBkieOm+M+CeAmqj01e+jOe
IGC79jSGEqOc6SVUHW5RVU8ybcsSQeNlduRH+M4EfOSbRCMlGRUdlkEpM60nx5HHNq4h8eDCxd5/
NOQ+EV2Wo3vrN99jRsZhtOV1i2yjW7rdJUl2bryv2AEemoDbi29MtgXBevQH/6GvTc/0GJsiwrmi
uomLMTp4VQ1QEORiR8Bq1XFX0XCvWlQwWNuH3VyGjYdsDSuHhNGHP90FsMiIVj/wQOLOvmcN9krO
RHt+vl0CPCDEJHBVw9pq9XvQvoYNUu6L6IIVnYGMzfZkZxdyzjezC6lv6vKwV5tDdh4yON7+guI5
G8LCgbl/+Dh95gvhX0QMbJ4TzL0TvaG39x9U/98ioV38aho+UyquKthnW6N0OIUENEN6L7tcOrlv
GEHEi+/wYwqWbVIgqwhrphN/DQmgNFdtFs5MlfkFpaVXlX/ZsbPjwRFr7Rw9OdAOwnKhO60/qPjv
Tpk1R7sKvpH5WSz1V4MOqpDwDTTflwkNB2TMHNtfEiRsMku9spSaLLuRIdjNiqjM6QWwYKuhIny8
mXrN94hbEZPsxMlDuqqL+75nQg+RPmULW4SKsQSf5iGlWe8s1VCUJyv8V4YkkDFjICQwMgnVdeFg
p+qyCuVI+UWWBqJJFQYxahtTtbPFisfXzpVhTaujW+MSw2izSTgzGy8rBmwJRJlptuxQ2l0CT8j3
DprXPBoIZmCbL+dPMUaBQouTjfX+LkRbER0WzZ0jR1GmjRDj+HdkXT7pOub9S/9SZNnlpve36ynH
PO87wqSCrDCJMTigjiIJDikPG80hkvYVe40TinHQLD02RwVPvXBBJuZsQLKZN6FCmeGZDJj8OUTV
0tAeuCqitbC9ALV6XYaud+Jn6aa0N/9uvoKzw/S9ywcl1nmuE18VzBZkABOgDzYI9g2qMNwGpUNY
4gN8117G5yGBIMCHWGmFxp8SP/FLAc99TPplBAqU/hYLhvHYtlpSvGM7qvViiEhn0SOeGgRh/UsF
LJ7g9m+G98QX+SUEYiKr+IS+wzDENakBcYjZqhCjca+h7TiJfElTgrfhIDzyeOm0fQxOr11ibKOc
/KRTS6DUpyUUgOM4buF7Mi3iQPkIzmB6sWj7iaIHRuDJt+QVy3SI1LJigzDcuNzyySuguqht5hyv
zUMbXVSYA0Gpdn/WjHhYKWRtpELEC4V+wJfSa9dzHMr3QHkFdvDCUvem2Z2NULxlg9euQH2mtymb
+FcK9wRI/Wo8f5KJok7PVIjvrGh4ygiHWFlsexLF5Xp//K2meXpoHCpIHW9jYb92pinAR9M7a6Mm
GKvuBWJO1QSJcSc/5s5hSeN9nQEgweCqH5OHPlJSG0tfW9zL75hmnCBMVvbgSbUsh1s5P35Vdpyo
x28A9b0yUW7B857rOCkXNab67yeqF6FgANgA46ThreaDoj/KPdAeB0zghrlfQSKPH3V2UcdSm8zR
RAAdSOpAF+m8uyB4zmYzyXzwNXhyKIM4MfY3t0etmN7It9/bp3Qp9piUZGWmnun2ui/Mv0PBvGJ9
uStYLKLmckdiVhAd+xovBnHMol9ihrSTn8kT8X/ZpasuwMCkBYSHAAq03eTvJctrD+hOmq64ZuzV
dc4Q2RUqX6M1WAETmIYs43dJGIBqSpOBpTBo7bBgyTpRkiVZ807u6/wOBQnossY68FFkNBt4pIJ8
Tnz6+jIR/19uHTbu0toCubtIXxYziOTrYOUGEwh+PG0nGpNW+JMsjfK0kcLU4Wv/ROZssE0GHl+P
6nHOTlzT74LoJzaT/fBsiCWw1jfhFHHgMa9LADng4Ho/x5nCZqylolIYtdd9gVR9hEbX3uiVhSNv
Ih4r/J2leEodXW5UBAWfjfKp6fV1AmhAf/n9XxczxCn12YBIqp1qI3X/6DImymW8HDDHGlGDNUWH
L64T1QCkrG98HI6VerVawMD6pQ7I8lMmTxud0+w/7SJjGQ1GEnjy/PoWJMafMdSp5x/PbUa3uEjY
eVODmDj/dDJVN3MRrbzZgeqBO07whh4GMBzAHM5T7MJggSH4BlwlGHaSkvCXmlL0EXhy+obzvTPp
fc5GHB9i+F+x7eoF7aSJD+zjG3vGlfSVIdzyBe1Y1gIukoQXXrafMyCz3rN+32ngLVuUCM52cfcO
8f+98S8+D/B4Jd84tvyb3O2PKp2I0YBM/pJRRAPz5x0rTmRdiZjIwcWC+81Fn2O8XM6zxXGI8AD+
xqPr7i1+afZ7T4a70CvHmxEpQDOWIwgFDaWR1AL/To2czF6b7CUgWdbb/WJM7QY1yXZdvJUbxis+
XHgpNn/zhUZKi74wtrxA1zUwRxvTt/IGIDfwTSUgb3D80LnM6Zae37wFx/AYLdKw7F+wDYcgDESz
WHOUVteynXtPJIq5aQdbhBG6CpRMp8Niaz+zIZu2woH6PEG/nFEwB17nHMb+C4+aV6EGhHv7LnXq
HjP5kY2MPKCJd+RJVozDyG6LUOmujMz3etO+AlYCqNUDElRV+pDS447aXFWF8CdICrh391PA78NI
cih3NBxNuAoaAYLHxoYsDQGDSI38oB/4ylDOwbH8ZHHhO0twchGtxONZwZK2TJ3urgj8+IMEXoZq
IoNA0b4LZ0Ho6WaHP/LiRy134uaB6nAvWZrQFE+E8tlUT02gva4QL6nDhRMJGUSXx7gjtOy5PYm3
IVyHw0MJG009AggFfkzTs4dM2w/U7smE1TDsymoMtDT1b7wlKPOqCForaN73M5Sg7wruuArCcRXa
MX5YpfFfMg91C4YncOCVQ33b9qFK7/d04t1Aqc+lK68KtLi1yz2y4eBAugcBkyJXjr1jnk3UtdV0
lnlk+RrCrFm3758PF0ARvB8hMYE01jJoS/NjHmRTtbr/TkQbK6Qih0+Dcq59xH9LBb2/Cdp4dG9w
vnDNSU7Xa+KV+WTUnBDz7tbNIVJe/0PVMTBJ21YGKuwf3FwfxkTxwbivTj4duMCVJXefRE0XFywI
M+gTKgWcYTopR4u++0QqsNhqGqm3qzu+FzaGycSB3Hbr2WtBftjho/yDpDvsps2G4MCs+JwZ9gTW
HxY0VWhXxy3ljlNqGj8QdaUYrc1yTp3+LYYIxM9f0tBd/Oqas86HwP2koyp8MAXKizdw0pBlolc5
P5kBuC+wzIoYpR9XDfNYwnuKMPTZZR3Ci07xQ8eNyDchFrbvgZBWsrlx3JPv2eCa2ktGt1HSmQsD
vczvEhxxZcYUKiiU5CMomNiPE5sAXuikfEaIaHdd1AHnwmjFXv2/PTUIPCA531jasc+Yt9bnjXXW
RahSj5HMQSE/GbjUCffx2bB79C3Dpi0Om+RUzpyhsDTPOzs3Yv7oAys7GcUCF8dkAahTVFkgCvEC
hjmYT+9LGmttrxcAeoLrTCmKeCnn1LPZbq5jKf0YfhfR/0RkoKmb97CdVW8yj+SVwTILgDz/O8nI
Cnxb8zl0MtI4ju6LpbcnkfNIAFK40rVf8SrnFYN0bUEPncvtOXSNV+XnBd2U/ggXQlY1pUbpke5A
uzUjg4vGqza4LlRd12dmgO9V/po4DI/tjCySV2sSDbSZtENnTb/iBNLYd/XS1tm1ghL9R3K9DusW
Mo/3E1fZbvywgVntkZpl3DVnRAavVlpvWPxlo/iKp5r/yyjsSBga9Qfar1cd+8YkAyiqdMYhH5mR
9yQdfc2KAJv+1U/PSaoOPLkMwlF9+dBLnDLfHcOuey/rkZB2Oj4k8TSqR/Uh+zGbhus9rDLhTE8e
1wjxbalazDsA1uqIKSGsjhA9C2gKXiihuDzFKlDaGU8wr2fzuD5CvZflCEH7UtCfat+PcVzBZg9y
kK9JhxQaC+zz+1RcuIKSolPMLIUFAGb1/kzVonVKeTsXtDZsxPSa/4acg7k0aJjgniIoHWTAn0R8
VnecqiY3cZLUVO1Z2Qm5Qyb67sSvVKyPU7dGP1VdlA55gZ4YO2cqjmDdBJU8+XmAgn4lNA01uYH+
fOeY0gmsHWaHMygCO0Xcq+1YdhGaK1bepciuxLbnp5yY+gTfL9Ba9naY4Tf0SrA0nhIxHdSM0nw0
+W0gdUP0CC72GT7WbjBJ8V01HHwonB7EGQqj1bZ2/zUkhR/JYi8rxqbZFuL6nD9MayKx2eSNKyQe
8G8+pmO1zwMLInikq7DiG5D3/mpbxkGBX6bAvWuPPLEsqiVYRF9NGm5moYLvlH+v0dM4V+gpYu9Z
mRkZAIWmCftJ3N+1AuFIEoNl2jbb//lnorIYKlykfACCkyHM876/f/uLHnuDl3q+aE+YzX51qkc8
M24q+pmquV5CBQPQEuqFAzxldekTqV4cjhVs/T4n2pbbHx4Caedvnu2JjR3b21By4leOQs9I2vsG
vafYn9Ue0ilfeceqUfuyYMc6bP2emebKAeuAmXS5DkS6DhlpRny+jtUuoPmVgHeqUsttHuDiTZWP
W3OkYgabI/35wVrZzg20SsJIMa1NRGi6kpzbMLGEpmbOGtK4iFhcTKlKHRtITk1FOzyClUGi1i6+
npiqOvzWoNXmgVhyQUSIOBPSnZwlDqCdnTku5dX/ibVMdJpL+WGV2B4xdepUYrTOL3IrX4mJJo8N
MilE3kkXrRtivmE//86t5roaxnpdIpEaB2V9+WFYs0nWvBoITE8kSW+yMTCPE0kOCNLKx+xjOVVH
6aGz99rpWe79oxtr3WC5sADnoz517bu/tLkTA1Qw+IacjFgNj7xxUa8SGC54DArxUAI3SrP2vw9L
mj9ClE6Dhd1hoP6/RNAdYILKCJPKNq5Iw200oUcRwxatOEAIf9dcoTyyj/5wVYRODYnrQxmIkOI1
ZF7uFdC/B/+X/9DN2CUFGYJgZ3k0kf97DLlA/YDlKTiw0p4gUWgbxSxjOnTz5Pn97USHQOS0RLt1
23XUcPM7D0WSc4elZjNb21XBhQNy837EnCNKLukkUnmf/PyHxOcNUtvy8INJNhR57RT3dPr/Ceb6
y0kxSgwAbn1sPKyO6UuYbzT+nfz6sbVXikua5zvzpew3OXosHNOFtGjid34NR7Zqd5zktC4SsTnC
fldK2mjuSQ82FzZ3zNOu4TpWadg/CMGiFs/aSGEMfHD4QOaBPeNnXWgMXVekKyQVfI7rZd+DmaXv
ryMdo0I/+0+J3Qy3XsLDaG2XKj8iDEGoY9RrNlUO/shdx1wY10tVovDPA0P50swqlTYRE2ri0eku
HXW7bbhScL7qu41ITgf8jb8AL2dcMSitS+huQT4Q/9mlLvREB/SIkPe6otFeDO2EHi6OZYpVAKGk
7ccb7IHyB1GkpKoUJINRb22vVxYqglCz8j5IPh+qzGXMPFQQ7eH4X17MJjNOy7fCXYaxoguYzvNS
BkB7T1/mCFPj09RfoYbSaqarBDXRP/bee5FNrtte0Klj/Ycteszm5RD4aAhMorYHPRGd/rl1NtwC
01rrfPzMaeYWcDIJdnQWvKybjAMxqdAIC8+ZqLjBCIpE5E3aKdyLo1D7vLvrC4glTd5UseyHapCq
QoeUCjs4kVKAp5RCiXBOSAWbPJGTSwX/Av8rDjAY7dqqIZ4/W72kBOlgoo9cn90F8bUQvNTExrUw
sujPIvfxpmow/nbD44f14/D4IdmFKgOUWke15zF+TO+/AWhFrxXOHgiVakQaAtzmjz0Awk1n6Miw
b/0Gx3DxCoh0EPpNpUN9/BObQK0JofljVFyp+HtJ4lMcDNVx5tzqNaokhZiC3gYheZxwOAhgN+If
4I8QPARPi8zbJHrN6Cz4nKZOUZFDEWYmBbToLuJXGnmCSuyA17aqw70UccW+YRHiTZQ+k3kE3zZW
CNPA6PA0V41M1xRbv1mzlMmcfeLtyfTavvJc1Cm8u+i2DNIj4NZTXuxCroDc4ao0q+I/Q1zRvj3M
i4/rwpI2PQANBG2UmeRvr8UEYUGoy1ltTYsQXlZ8XexuM9i1eifke/AQD191Xwts9dXtf02U2XCV
ZD2GDt5oOd0bW13GwmF2p7wTIcZjTPKGc8hBpP+tkKDw6haC8r/A00XUYyn5N4dAS5lqiEjgaujY
lQjADEp/EHYu7UwPA6eu3Ki+iwp7NDgeQJuZPBrGHqqDR8wu9usJjWw+FrDmIruV6yGC5jKMkEJx
rzCyvJ5SuHeR8330SS44vuLG4Snw8eMPctFD2HqqAo4sJbWY9k54So2rHiRA8jrucWU+GDdFi0bs
+y4i+VlsuEdB+ocon6SZFGKj1vjJ1Y5/M2XlgzPyfObsjqf+J0cvAyv4KzwL/l8zUunZZ+D69IvX
81g4Hu9ukdzGmMlHYMby/gUPeX7HnHbD0Gr8PRy9Ytpu1n/xP9pltHWroJDbHx12suM7gmyEt4Pe
Yl/yYfFy88MoaiVTYeC3JbmdQD7egy8nAeZxrJGCxYW8jsUZgIhCTccE3MJv7B5hGof78VrDmnIc
4U7imye0+DH0rVJmfBhwwAG3IUBnrWtC0jvRdu2o+PPjRLN1S7eq1dw64+rLa2KS/ltOz10ojzr+
/kQj8hrVz7IKRLlcCw2iUBFm1DE7jpl0QVKotT4FKtVKKZRxikhFxqMPbq/6fa4jqbfJVc94WPKJ
MeAQ/YIwCC81iERfvX0/1n3G6+z4R44508HWXAbq+h7ICdqhyqFZAba8XneHvhJchCi7XPkxqYOR
qYasIM6mmhSi/BwNAX78h8I1DD4AoWXDGSZZFQ2EfGyMGx01mpTCXfi8vKlnNB5537iJ6pHp7B55
1eP9+40stjsY+1Ql/C6BkHvD6wnvkEN90GkBJFqeUo6stKkTkw8rEFdzshBJe8mY8TLgPtybGO/A
L+H1474SCNv9lTgx2sUyzpPuSuqIECNZ/P1YxKWiRth8hQMElkkS/dDvdAva4m62DKqWJo2N7nLV
WUc8PGsgcsnyEuJitJ5cPqhzBq8mKWlstTKBEXSMo5b2k+lJ/on8ejeFLPbtY3YUDRwp2NWZ49Br
xIhwYvATHd7010FrWatEB0B+PXQ7Tkjcu3ZRUt2DtXRS+zyz4f9NPGipM75FPMyQUqQIff0xJiS6
IdMo0OACOr7XRO7jpoQ04KNjQbTKUd9qcYpneAj1Gepy5ByNzlrdSibfmHy5twm+crAcud3czpYa
Tx3D455pn+XCsg6CZRbzTV4h+fcQhVffqS8cV2XomnVA7UvwipF9xwOi+mST+8Dv5dVRX8sJjdWu
nwmC5DN01GB09uxGs23lZ+g7T0v74OXOCf09AIlOa047zQEc5UrTF3AfnuK7CGcSCo8kC/Ae4UyD
k4+daQKMQuOZtTaMsGAmvt0kW5hTEzv10rzI/Hxswe4KA6CY8FCX0nyqBxqXa8AoofjtJX1rl3cJ
ZjB1l4SctqW5TVRfHUlWOrv4NJz9iPhv43DZFWXETqVz82b+KU1Uy8lX95MMT4Cgt4U+Bn0S6kIX
x6LoYcFiVtxJ9AnbhB6hGfSjgM8VFuY54G+v9DMDHiIgBUaXMjt9dhlGQzY/k/iQUrFTBwvJzZMo
UpjaZmMel5wtvvHedkejJHVdd4SmRbitVJpr2KdF4Oync3vBjOfJpY/lspqtQcQb+tnZh38JjrDW
1KdNLddYGa3fNqOmybzqnaXGfUv5Ro7+LIr1pjY184LWG1eYqTccCB5p0Lej89sTZnlw9p5Nd4OT
mDY4pjjhzjuCmN3IAkascpzlVfUDgiBuS854sdTYgU85RoUlJPAU9Issj3pKM9KWdJcKfzaeLpSk
7ZOo3L69D+1/GLJcSVlRmu+JLECaMqLWv3lFSDuZCg3uDjodYuhlJ10WaezEqIRjobEihCL0kLxt
0vDpEoUvVQTQGcu8zcLurNlPqyUbrHQagalffvMHlbOutAt0xIqjGnTzU6+ylUmeToPWokMZyKA7
/lVtmvTw3NIjLqxLkSSa8qv1z5j0qvx8ikmSNdbPYV5erY0lzwqjvKaa7dxWPhoS9qXGpahcUwMU
JrwEPgBjocLWzgeigwyTbpYSW5akJ+UpcAULPQvM3gEwrkiZ5ykZ0hVZXeBVKQC7cSRbdnA1QyRj
ftZ9YAZoJOgPDPBWeyiDO06gITEQrlp7ySVD7eYkmCJpY1QjUA97dXdE0IdpopMg+y2O3a2cK8Dk
fp4KToM2swPx1/hxCJv0VVC7alEAO9NU+g7P5DQDULQP5uEFSwNoi8gSY6xQnM4m9eprLrMulL7r
2t+s1OjwzcKHHkR81I3tJzTIuSRUv5ngVkxdwsg5jHktArUyLQxNyY1FjUPP2jSmKMExJDtseiZo
iBStbIoCJWnDprAE7REGgiUiJlVzWIcWyJI6qAtHEF5g8rzNat7rj6XVxASL1o4ShbT/jNalQIwG
vxhrXjGyXuOJ3hQrmvbj1hKk9xWHjBWMWOzrSQfZVBTzVPTEjEj+16wp2rF9yWaFJzsBMya+IcMo
ZEvGhGevGBtgUmZlchqXuMl6m4HFtzxO1E0JfIWTcEFdx9nr+WLdrpA+B09o2RW65sCz0x8Hqp/f
/62eNxXZQdXNyV4v0io6A1LtRja1KRdTHAQdsSkgpvjcODqLZRnueuSshnGj7KndKXua6GVyv7po
GhkpLamXmN1caEMR82lBrsWfN+Blf8Yw4fHSICu4Zpy3jwhwE2+ZTJE2HnVZoiYrNeIA0SZOreya
zihStlAnVW3fJOpT41egaKRSOln6om/JUypt3FBfN2CCfqltixoyIZQ6lG6JAMFS91RAVSbR/f5G
HKHYuHoTMF49CEyfXjrspo/CUVGMtb/tZlNFjnBipSnNnCvarORHGIiSWOWafg/SWtsj11CXagqA
a9zTnBVUfUeK3QYoJ7bHFZJ/HwRNccvUh4vWt1uTYcoMksOzYSYlI4mc2gMFRzSHbVpO7hjrlKp2
sjBDF81z2rlTDtpPWSnQsPk7+HmPKwVn44aRObo3UdSfoEQJYeIDnkAb/FTQpHJDeycRp4yRSuSq
ZZur6fsWkVQ3dpEVvkzk0Yv8yhEyr8z04GdyV/KxfwTijuh8nCKV5vhj1o6LE9C2jjDJeRlzBhIN
y/PQZbkTOgdnbdftySE6OeGUSR2CoIJLlnqIODfO+vDm+mCtne3hL7E6OrLnjE+TjBl1Ef/DMZMd
3Ef62Js2v8kU3352yplhPgiL63FNpOWYUbEtaCdCiVOV2xYQ6kWYQj+bjoxfmnQIxuuk20ieDhWr
cw7+CCIpUcPr45GLEQt98tYgd4d1+sWaXHPsYQGha6uKux4XXSl/o+WDrv7byaUxXBI7N56qZMk3
8iUgTAP9nyUWOnkaxMPcmpAjTbJFSPSIWtD5Zk6ZH9CrFGmt/R5XfjaAReilz3LYjX6z6PC+g6da
e5izdu+E8fcSmuDNJjtVeI1U/qrCKcRwzYorZXAqQ/9UACxQY6PgY3ve2K1MfRE4CVODpMXvzfN9
C71iflgCbEyxlTk/VZU89DuXIR8eCivdLCaoB2CsOYkRZ54aIDFz4EPj9n06dZFu7LWJFnntfEox
VL8WfLM0dWRG3lUoaumeijaRFw60QCFFWanFFSml14W86D53Cf4rKYwVFzDJlMm3RvjjdWPITPeP
xBqSQbQZeMpmjsVfMF7as9JDM5wwUDUY/kuAvQBIxx4sYx/wt01tOaEOylyEEfEkcah6T3I/1Lyy
tzOWFW2sBVaVG1d215AIqRjtHpf+w9DM/ZRfM0TvVOl1EvjIpW4auFuJ9a1ERhOxSiBErRtoc4mS
YwnK2l/N6N/vU4rVRcIRu7uuBoVUvEdo5T83RK+/6kEgpgp0LeboC9OSQhOPvlXOqWK/jDqcFBD7
zrSACMUx3U6qLo1ZFYUEiISUjudCe6roGq9M0yYnZejS6PAOPM0czVUxfLZHt2xsSbQ944/qi2IX
JJdl1Q4AUN0Nm45XzJRIVtLLkSHbWPYwrHLW8XXaiiClNaQLvwWBl8qHNHFq2V4ixuJZ6HKBVk5i
9hBxC7gDSizPQinMh/UCRRVHpTpbekRkSGSFVgEnRW3Kcn5JxQOOgNHTJQy8PhhInyH7h/WN5EkO
fQWyuFh6ODnWayOZeK+Ym6hx8orr5AGYN5XrsgEjfWtaHz0Myq+5TI+JrsRobIBGKKwYja54cvnx
pcC4e3U3JkU2SqZ3D6Nj6FNpAblSeZgUqP3XPUOOVUxGy3KgLlLvSEA59b6NQgOiwsF+4JV7CJjw
SdMep/ecKo7gFhQCFYlAfype22YUDdNup8cbBZFJkhG45NsEoGd+YCHd3XXexPJII0UZFuSKmkpJ
dA+zUaW72FYvQu+D5lCEVdusUuWeoW5Kko5xm+zIcGIY+p9RGq/p1/IepsqLyy/asy0YpGSeeyyn
KW4a1fjswJCIo3caxFGrr66Cb85tCt6T+noRCL5vMA8F7vgh/VXaDN6YUv5L8/Tp9TiFD5agdmos
N7ZQLK4X8h3EusoVTHWSmo27Cl6y8xDBRMcHA3WIzibrGX38E9YHszTRkQCgRuF/kzd+ijhm9uqx
pxQYHMG3ZHPQlMqy+J/pSGpXSwNj/dVGxyYUdqRSZIyr6IzvG2HgdH0XyCtwhHcDAIzBPseKdI+x
nUQS+aBVAYnfDNTeGUQE0DD0vjkiM/TpPNZLyJMN017gXYMH+11CwnGJopZ6y3Qk0me23MlM9+5l
1QVQ9MPjh/A0ftYdp0lWTQTII3+BNpShWRz4VH3BaUXdzoi+K/GzJ6nLGjGOqRkMn3qYbzSo7XxZ
/KhHxQKM4aunzNVc4TE592+5S9/iLSmu6OR8QenrMhaV3JEYX9KLRVDzZESxJODtqZcKtEWDe5Vv
LzM/Q1H/fc4EUaLMvbcIyzKFDjJ8K2do/kAtlZGSwh2PmixGW8LNu+0vd4OZyaBucyrEgaa/q1El
HkdXT/BVxOfPtAphi2BJ85n2ojT1yLN2ZJq1VuNpC+2NX9ajhca18NU3SMfUpm1UFgSH81bSa/ip
PJPxw5+iM8gIgAlRknrypkttx4ABwZ6IfEwVn4MSueBI1rcxVGnoOCV9AiBpw7Oo40cQXA/COB8I
qEoNE/qqoulIo2oK4shqvXe+eqlYwntVjA293AbilVQKA66x8QutR0YTBQZaC5l3oe3XJML5jQJ2
/v5k9zLjbCMaIcyU6KAP/mtwyct1FkTrvhUJVSO6GUmmmFaSqJfJeP6ECBoWpozeBafqj+Zxhmhq
gZuarXLqBn1ic6AxMp+Xp/dKh2Ztt5EapUiut/2XGjEWPUv4InxOL9Ed5C18FQOjJGq6bI9bWTmS
jA4/ZPb4fZNJppjGw5t14rofxTPesTA4wCpTcV46cYhpD9Pe52LXLr+IY1TdYL+sk+Ol9opeLXH3
SXHN/vmM/F9FxJWhNPpkfy/2vIvenQ+gLzX0OCFcuzBjEX2UOu9hX5siC6VT5jgS9i0M1FE9YNo/
RRYoz04nEk1O8cU6ZRU04vdiyI8C1OzUGsXf/gfKR+rhemVNMyC85vyyNPT+WJqVPGtGLoGtdYOc
CU5q52HIgsKyabZjyVh4hM32LSZ9jxYZga6UJ2a606e0FsyUiLdCWXmbxFCl8rgLtSjjLL7q0PfC
W0R7rINAEEZuxOBDaxxAM/EGpuL5iFHSzIc6u+pQXwcr45fkYoRZ58EopFEqm+ys/URdZ+9+Uqnv
/cYB3ndhlPcxpxDEvYM3V4PVztICSmYKeiA5x7SD6RN2IX4uw6giDxP6GgdvCRPddHv4SBZKeyjh
Aa9eKGTTgB3Fd5lw3OlKWX6/d5yK9usdu6pganLuerlIOS8qnT996UCa2XzSLFAm4p4saibemBsh
sFxUWbcdEVu2R5110wIvKCsSrEsmZhUnwVyljT0w3Egxrutkblc4GWxeOd+QvHtUOxZJw3sLNYoV
yTduzwTahzeuIU5fb+gt8WE6lKraJMoL3Z9VTuZhUTLaLQQ9P5bSi0wSc72zz6ixLLtMmdPNXWq+
6vlpx/gGDt2pxLDZr0dqfnm4PCcmyv0aUHKw55e7BZi//SY5nuBU4tM9VynL20ZngLPPiWoQYs6i
R2yawGIH/p6khMOdCAxkT9KbWeP5byh+e6bymHOf67qydH00Ts20/T2V8r0hqrlYrQh9lx8j5rri
m9gEAq1xwcS7A8L/Bhe6HPW5qwbHiPpGPwdhgfdquF6ArIthvRJtbctis8Z8brlH2D0Xz7hCecHz
KvvakRtPjBGFcWut2o8/1y5+oX++XbtAvipEeOCEKblfIr9IkEPecxWRolF7MF47abE9ZV42Ml8O
pJBqW4+4izuUjI1+HnQjWQcuWLumCek//eHe1c8bqZcupAVNFjD50m7dfhFPZmRhw7IqO2qZ2pYW
7mHQ3Ol7NVew043oWfUjvGmj7I9oOK0ueAL0yjeb0QW+Y1ne5XJHUPLBKzL8MsXtBDdupU+BK3/T
37RGGwVOsBMznCZIYtaQFdCBVj6PiMoWCjoVhOQeJ7IFvhCBZYqLam2X2iBRCwO3NsijTkV+b/f5
GCG0rGDgjKmW7oO0mlCNfD1PvJ+xRHjXsTewZuFrhpkw9JAl2zoWHDcCOUh8DFtMT0taPm8I43uK
y54uCS7byLNn4n1hcdJ6noR0SLTNh8vmTwzMrcPsBUmvL6IYhWKCbH+7ycM0ZXZYnBSpksd9B/pe
Tl6Nw6AqeHmwNVCvhD7TcAXA85XfpcVrHY2fdLqwBS/eVzdKSUZMI2P9h+hhrok7b56kbJeQSOhE
OGf7OkbZEIhkWxRgAbpLgaoDUCqMQfQDJgH6YGUAdH2RX3+3gqz2UATt3px5Pf/vpbtiYKpWGdrs
HQSCgcXWKWSLyjbXjdgNyh2depXu7LAIwPLhBzsM4go6Qd/ElW2KueAocJq6jRxq/ZzrnjsCIryX
/BfYuGinLbYGzceuLMVlYms31P0N95llfv0dAXdIWEiPHsfXLnrJRPEt/k+ww60vXGcMSa+/Cx88
C6XQ0lsuILF/kvKBjSM5nAPx9/FC30cI/SbkBh2APtQVYtFNaF8q1CEgmpYWFNOMYMon7LP4T/L3
Y9ylkQADnh8L6Vna1uLN6Hw2pZBRl7TrfuXsw7hM8uhekUtNBQxX2wGBpaE9WAXdBhEN1iP5DX/8
NygBZTX5KF75XKa/7sCCU7O+3CA0RipWUcRa5+dQSKpn/YIyqSO/h19SD+8EpjNapuBEJwlff8o/
O/+k5hplR5qgmi3OWQSbgXe16dMTiH4F07inNeWuTt5Mu1eVW+tIpUE4swHsizTDRZV59qwtOD0s
r6ruoKgtf+lI0DmFOhApGY7BacDgqoNVJwJ+dhxT53DrA0r1aYTQ647NwwTKhALnJJGb+/UQUR09
qKzuZ+N5NxM7YbOBBvBKyzKCaWugJ2g7CY9hfwHklk7gzF4TEtWfp8txwy4n1k4s2Y+xoj3WZWNQ
uWsRUmRtQtiXaLM3BiPWH0430CXDMtSmcn4NadrOJw7dkX9S8lEhiuWWffhCualZs0DZp+zwO0/y
QWG2G0K85YDWRNG5Ds1rWC+mxJeqVqxNqVX7sDtngqzj44jQXIiYE2bW4O0SePpTGKEqqvRsBEWK
17XHUVxHwHswVblGwVP2Ym7ykfXJ6cFD3A0y+Bh9D0IQsXFUHXdCm0Updf2azCWqK750KbmEXKVb
JrnS1/iP2MGwnKye5RZlr85mooRZFQbJecZvKUTrO3HhZv92XPeWZX9hS1zrz976BPzYvErGgYuN
jqMPvDxRrP5WEQa+yvFPYjE0v2vhTK0l3z4flCh4nSeV/Oa96oM7otkMUeW1NY/i+9UgNClEfgLr
686xVBYrIqNIssIBN1fLp7oqMy5RNbRFmoStHJJk2XCtY9cUgZ/Lkl/zsnIpMF8X7h6Dumc8G6NV
KxW9OZMuv4Qvpgvw0TiBF/3RQR7XTZaEnbFHD/xqRSjGk6M+fUL2HyZkvi7D87mxi1RcH3yVW61+
mOtQJZoTDkItxwqgmUmOJ5zI5R2sbn3eeF1U/x1dbwnnPEGwbiBYkaaB83cZZxBVBblJflSQOJhc
8ZFBxvTFPd/JkQ5EbR+yE91YpAC4RRQGIUunSUFwd8s6ai6XDJXGFTvbcbxB2JYIH+enHLiDnvIA
bMMhp/u03JHALQhKnoMopwkaLLR8iBLLC6jLHWVUG00VPkBuUySq/mDm91Lamn/YsOms9EaRN+nE
oBdRHEVSogBTqdZgDb8K4s/Jn9uEG7eeDVxNkIhSvAlQhsR1AbH9DYokUQIw/Qu98LE1Ybb8Rb9s
W7SgCwPQfU9fFXcKH8YaAuhGA38rBN8lAaJlkFdic8scc4ZvTbCgWdi2jr/HofTHelnc5F+/jSVY
D5g5JDiNRDINFiCxHeiWhBUJbNOVz7Kqs+9VfeKGKZ8mPTt8IvLByjk2rEWlQevyna2A7TZoOdth
igSOMBkx/7ZGXwE+RdyttwquBLZxp2FMDprvwAz/S/9wfwXJIeYJThF/tf4QYTKwT/DqTeA2tbax
QPo7oySsFT/S7UcIQbrBRnzeBTUoZtX50YyfpCWnFn+uTcFE1X1xH5YHuesA7t5hzOj3rtEcQ6kZ
gPFU2SrmFtaWN0EQQiTgY8w8XlffzHU14UYYEosGPcBXGb1QQZCRejKgc3lIX42FgQc2jvkpc4IB
KM8Ns8Nee6/sn/LyjmeR4ClkMUUNcWqUCFNc0v9/mZDSl18wGtJ/SVW+2TQpsTMrKVEPp5BHYYd5
fI29YLvJg+cC13+cP4YQDX4QCGLJegF1oQ/gUrqCNHoef4r6TAFfeydthYtMYGW8BPBStOO4zHrn
1k+bbQoxYdA9UrlN68hAXvtiyZeXaZkTsGNLBbK/KqmwLqO8YYECuDaSQmMEHORwGXgLUNEkDjhg
wYVVUlTlAWfCvkBUvvCJFCJkAAjVaQhEHivSZmLn3Yli2P8tDsmGgJ2psZjjqbJGMiG3I0z/mjlF
Jiji2P2BuGdrjhMpLHVXXBnBPyx8vindEyYScj6kLWEaeFelEyIQ/oF+1PKCPW9eSN9nHQHpFtyh
J84/7QEj3OfHWy5ypS2Ua6kjemnjuvFwJnBWH0RFmFI0+Lpvk/kPD2dZhdit/i2lvx42MT7zl1Ye
DDOMM7YICdqse3o4SxlG/6+JQeiqQ8GLe1uQw1Q5eDA7ZnH0ZNfRRgR4QA00uk4UWczgpISxtxvG
G40NNE/h24JeLIrGZAbYL0uN/mOEUrZDqvhPD/KAMUcln5ERwnoaw+pe+uHcK+/txdmxNPUCr4bL
ifgOiVLAoACRaqUMdEJIZ3eNlCCLCIC2VZvUn2hAIyloF39a7LtIOszScHXJCiQqUs9utE7Rjvga
LzmatIrUkDjrMA1O8gYHmOCMbKPfKYcF48Qb0KUN6RrfQkQ6HY75mOf2yPo/l3afSfH5AaoGz7BI
Cn672g5rWe3YjONLpEBzCxmokfVuwJ8e8PsjXcGnU+MW1PxjWNgB3Elr26hhFWvjMnXVt1jrK0vw
4fV4qWl9MPg7vXkcC2G4CGsZfuA9Ln8uZjtzUFtrNpyISYthgUUq/RBspLEEVr3aD6qIfynSPKMQ
jQkel+EIUgS0y5kp/o/u2/VjjXmvysjmVzsuTAS7mPv5ysH7oM60qtGVSOmnpz5LvzEt8l2+TN/a
msxpdGp/HPjsHpfbUxMLiukyX0EcFN0pFodP2gH898gn0u8+AWTk1cm3fRPzGSW05RljcTtd8gW3
WAJUw96umWs/OdhdVWhpV+7VaIDzVVA/s89UXe+SNGvwXNocnWkQgJqI16oLdhgoBhVs4HAHQdGs
an7iIikAKw4BLumCc0Of9sPPq2+rZJxjuvIL4Z5LrnLWcliW366veNCU91N4U6scPjlUo8Z8YUwr
M2nkfiybBQllJwi+SxjX2XDML+sqwaqERCcbAZNEYGpj5D+Wii2l/tTVRPOZEAuvFA2HuZZtx5Eq
HXuutCPPPVx/GvTRScQM/+8b+A4xIO26pfOG4SQos7c3AJ1Gntpwv92tYWAcHeTHk1e5+3olTtzR
u89+Ip02Y3E1TjR6UW5hyUjCsgKNZII852N0rHpm6/hwjAB9GNgcxwvqbveMB6csqfEBh429QEVK
3FzJDTJn1pcG8BrYliBt919PmGtt2AOQzvHsJ2Egf28rqQdPXi09xWby/jd9+tHC9vqH96hGho1H
pZ7LUu2Y8p4tjDgiNjscXzonLcIq/OrzC5NOntBOWiBvsELee8g/U3K2mvJEA/yvsIl8mrirgbu6
YlQiV/ip1McUYvgyD7QR45TqX/2qLc926SzGmsiWP8OrsD7i2mZbRx9KX7gBotZfVOIQ80sSzEUr
d6C1RZkNbOlKSAdGc6rOAYrBFR84sabN6+331sku3NvBRLSKTw03tPQ8wdVmoedeTxBUw3atZzDw
uuPE30dV/dolSLAQ2IzpEf8Dfh+9t+HTouo0+guCOq4rqkz01BVPJiaS7Zk2l3hibNbz6B5tdAdh
v5iy0y6/Cme8x7Mkw1C2hS14pO74W2s8ZB0IKc8pyS3l9PxGyYqnd3Xz2uWDFTrQzCuy54zG703+
5PeguKx/ZbAH8WJaE6mN11U6krIHQLHill7nKrC8TVYp48GR/SGFqo0gcnuIZP+Au0S/QbBbfFob
4iRklculdsXc1AyItUK0T5/6jnaKTSrB/PIq24PayZWFuJ42+H377sQPhuGWNU2074kVu3zTB+Ag
D3uhDOtgJ+yUMBYlz9q3UWDspFsEWE0GhdzCUQjs7CmDq+nfrjPG6iWEfa0UUhOXN0FRx0ZCY2Pk
GHHxdTV6i0RAaRn4zhKVeTnf7aItSmSLeINle5SnRmjwpSQJ1nzVWlgpcf30EbEOXCzMp31wSGww
hzIj1J6EgQbdvm8KmM8YSXMYDdd1gxyQ+Aq6cYPqJQaWb+/IRyZymicntWcb3fs4rtiyjB2NP7dK
wr+Fp7SKLdv/ayp8tOQn1mMN/hwAPwCsThnFKIfLtnVxLD/yNvb0tPB9yAIkSaQzh/SDaUUSuyh8
ZggnZA7aksPU4J4qhspa4UMCPAabo2mPyYqq/JjEn35c7fE9URmHQTmq8CwY/Wt0vJ1kG+zjpJbL
H8if0C5wKUKvD21qcsrNHrxLeHpDHxcz3GE0ecHtTxiyZdF3krJdhsZLomE+e+Ta5YCDqMNbSvk3
wWgDzYAzBnKaAUddx27viDcLlDsLYwNgMCqDAaa2/gOWhyvqJZALwvgEG9XWpbv85KVO2tQJbZE9
4aoOMVunHlGfKATk3SyHUzdSMoMXEcQxpBFZLbfMkwIWZbnw1MKPu6ss5XW9+89uLWe4VCfO+PvJ
mBqWLoaSITylxiehdY/sCxy93QtOoyfSlbtTd2NQ5pWnAXSB7+wzjPdfjFDS1y++NMXVuUX6XWzD
hWwywZQd2ZoykzYjxX1ujHqU0LJs16WJ50ePIX97+Pil36ug0B7ArZUih+GZWcRbVqk6E5Q/yDN0
EOZMfHQAyA1uFyfQppdSARcc2V+1sIvydxWLiJhH6FjmA/cmKOL0tEhgCpQILbSnSk2oNnCo/kab
LGSLKcq8RiDeOEifWDcPIQRuJkUni49ANiOFq7lQBsFTd8gJNQ4k1bpf40JpRUArevm3iet/aCIe
okMLnuJ4gLCKLsZjgVAl3V+cL6HTsFIDgnLnEz3I9tkg2CDI+tUXRxu4v9Nmyqk1mTpe/vDI6d8z
yy/EfzoIEPRcNpyKNGmKFTA08C5KjB49M3DIcw18NOlMfB7qFGiU/53AYCyT9veyeQ9e3au9Nvxo
GtzfXlogc+l4THYv3xcHGOTNw++UJqZJd/jwOuEee5L/QH73Hm0JA8Adk8XRTe8Tx+56OuplB+vx
IZGTDSHCb77fYr4HFONWflH+VbM0zYuA6lwyBkIR28Gob6G6B5t+4EM7G5SLgojIEqJ9q7BPr+7Q
xwLe6mDLeI9wH3oOq+illbTbhHD0HGiddLg+EqHZZeQZaaTwsmLHGc2U9FIoC4Qqkl00bDGOz/BY
VuxXGoaUoZaUqZcpKftXZfMYrEkiLL6dpE0zSJ87oFFEBFA4dbJT455/IAHf4JF3LirMC3+2upcs
iNYafXGoG2YqAmyUUze1wkVKvBjG7JbHI2+VZjZIxdkZ9/3qfD6IauBAQGcLHXlXdi2vj9LrxTLQ
DlhOoPkiuYGrw2qALjmNatO7WMuLOnIeW10TIPiDu6wpolnsMrldAqWDYb6ddF6Yrk9naQb5Sxoz
Kk7T0cAK0lJdGv/3WG/hg3P40Z3xl/CBysni0JNvGhquLKSs31mUrVZgMpi4oOOIi8n50yiEMtRW
nSZIu8ZjwQaGO52+EPxAH2r/hpK7BAmiSKiGJrh33egGM/r5HiPXwyiAi2If19ZxSMiwfWFJ5o9r
tVXH91Jg22xiof5X8diaVzGVBku5HaHItlNlAzmvhpjYD594uYievSxskQEVDyh7w0n9EV90FXgx
cr0qoi4UdyK4v8FJ5gPjVINpYy4vc2YLcw6hkT9OGWqugnB9aILwFF2iqwR/wTgbfwQbcvhl3R1s
WhsrACuPMudMwmwh1dOW8IrzhMg7/ShIVceIoaSne33GvQVDtuAHhkmHzcNuGCkmzvZUlksGwNtA
W8jZuopQMAHsD78bz7dhmyKbaRXGTLhjyUXnlP2EtdGGNJ1M3b23MDub16pH5p4CMgZXxriMqgBm
2/0SAfRk7ntcCPrhxr+MA20bCPHwZ0yRxPydwsBnuV24+UKp5DwT+KMcGSOASJza0u0QSuPSHMPO
+9uzFjiUD30Dmaru2sw1MsGR2M8u09gYaVAUyChMpZsH0zGnvWGXG6DnOQKwRS+68K6DkS8KBJOW
TtLwtyzT91xRP0HwbdixppcEOZ9ALyOmxK/yOdFFvduqn9EPWHiAWlXYe1jnc6skiVbnHEIgeca9
DNptRXu1hdZyo+rbPzYAF7VJVSxpp+PjbwMtvoGu4z9AmyNiF1sItMuZ9jebOayseBAe8ixQVL4C
7lB7I3a/sTfxqt8u+Be6UED1yqKlenMwKof23Rm4HTUcH/heTAlhlEfPzKxhXyxCbdTxwPO8LRuJ
ym27PjwNIK1PUTRh17t7bqcs6p+yl8C7J7F47zHTT3TJGQY4N23fnUrJbtHNSCCrHkRhPqNu+7o4
8T7CHZ2rTMNZ++MhX+2Vp3trjmFedVVQqBRZbLu40oDN6LqTYVXtsvRQ9JQExpn7sxyYT1Wygjf7
RsTuRKmnATuyEONQC1cs5a7pZI7yU/STAHAC9FilBzcTsGGwkz4wDI94WO0r+WK2h/tMx1CbolbO
oVd/8tu64YUDKkP+p3VFXP7W9XtVLqBov4YtzgXwNzyqiW4ayWbFJ7s4jSs0A+0nyL2Kf2JSf8hq
/QowmYqs7o3xGcmAGDV+IPDctyKaXqz32a06XtiMxfiefOteZLlOhd5e6MPHKkRfXtUlnRSV3z9+
yZut6atxiB5TTZZEZBpNEEM6uta8brdK7LD8tSgEI19qYP1M9blk4O06k/U0gkq/TVO3np1iqA7+
rXnszoAEHaPRQhf/TxKtj4a3hllZ/iMAN0Z5CfFpFQ4W16Kk5H658UEw34gXvfPm3avl0Bt/PnL9
BvU6LwBpDSfoN9oA6oFRxUr1qIo5LRzSpm7uWsESNFC5/Qw1m9uKf7nh/6LxO47xy/93d9YUPqfy
Empb/i7gV9swMP4n/d4W0TQJNVCJqc21R+Sjd7BTfqFy7gwia9LkJVMFl0dAzsm47VAOwIZ0GYeH
VCGoyXjaQekO83/JvpcRb3kpf9q18p/bPdsB+CHfK3K8GofKOkxLkUKuQhVhIVumFnzkr8aAvyJ9
LR8K9YQfoBcBgGk8Hdev7G+IvXxJ6hpsp8IYiTv3Zg2drCpYR8cun1ZvhTKYosQsV9lRAIEOmXgo
MA6J6CrExxb4vS9B3A4bouSD+kkp/sZ3MMNzEHwe5rVFU8EOjH4wzr1Je5Ac39qYrm8CPSotKItp
gSkcz40O44WTvqBgnDA3X3eVRRrRXaEmjINUjmwGGEGgjj8LF4E5/UV8qlgj2cx7MtxmdeZp6+W3
YCYGSqfxMczhW3jrPI/NA0YQinyCOZ2Eu6Gr0poj3+O77gBWVihrlZE8MHohwF4CTs+KGlxU8xhe
sY+fPf9R8jAhsVomC9w1ryNEKHrc4h0SJF6KJJOe0PS3W7Z0LMxBExatHEJAZ462Lg6T/HKM+2UM
AnI7DKh5pKWAPlIIKvywVQcIe5mZTk8pzSEns1iasizwGT1uoIvdxGYufc2A2lxsCSRoG2k6qbss
bAkepRO3lbtJTZv+RSox4ZiruKwySLUdrUQ5oIpKu/jeBq8f3zT28j/CvKkcuX7bc7n3VDjnR0/O
8MMfceDs/SBsMoMhqogWgtG6p6CkAvYty6j3zrITh/hXNP8R2l5xb2/o9AiwRxAY4x8l/pzFS/OE
BK4/lOhsnlWQpCDuXRw8gHtKzGgR85I3jW1V1qKpEQ1P9zMeBl25B1OhKqFjxAuuR08iosrvg40Y
jY5IGHkzWgUndk/72h5XDXkKByuHmS8XPTKyuB0VcNGMDYyFk/qjQOmDgbyPOLHKyH7hZBT1m475
rW0aRaoJ2GV6S32uKtZO6fseCja/7+F0FiKyszdYptkU+JGSLtHZxp1Uh8FMBMFAThLAtHSOQ/Gd
kNHnxoEKs1kvtMTtajS4/H5yjjqM86LPsY8UeOvtNEvv2KfltXfyPdqJ0oWkmdfdRtAUeylEZsLX
5ZNX4xDhQjfvKx1gfk9ZTbzPT2Fxb5YSYuFMLFx9lLqLnQAsYkG+ST8otH710mQkpUL9cKWCik+O
JsWPI6dUmAYPxO0m/JHzPn/igSzA+8wXj1vhq1oBOpAA8tOYKfQpvo4sf11xeLw6FokBgX54+I+D
7hVipkuD28eJgCmyr69o2HpS1kLz36LKmAov1SWQp4+uJTw9Op2Hbscd4xShS7KdEecl/tTO+3LK
gLdgkoDxVgWjXcoTv88P8gy+qsmsk2/Dxra+dP7sBqcJf9qPLOvZLV6L9uOSqNaZmH2THrpHAnDU
OymlDTzz9oTK0XIOjrlvYAhZk6RpEBs3NTYOkw19TnWXBdYRSlZ8hbF6UPEcmu452XhGJf+YLd6K
4++9nzjJnJv3jwbctM+DUxKas3zfUd4irl64VLvZECVP+JiL7rsiQI22cy260T6YNQjpYISMIbjT
4H4QPz2ZKR63eefgpZvMkL2qTvdcrNd+T2BjX2y8/wXh/Dw8dcBoXGBcaZw9h1AdLQZDcHjpg8Ti
stw/RyMHRwmmuxkPSWwOppTBvQwYMTWSkRANdakPFxPGW+HZo1s0j9CIKMCfgFhtlxpSHIqp98Vj
DBHwyMJ/WgtkG3LZPrvKUonrPOOR5T1uil34uHpl7p+e64CIn/8miQxG3Dz9tqu7HtOTSmH7KqmX
qCIfeafCT1LzgQJSkSWQvtFuP4ueK3aFJzUIyF97VPLOgBEpvuC5MtyMv2dz8YCM0/AkgVRwlgB+
vFuv+TdYf/s/Antgn7+jNlyFzd6pA00hmtwnMxnsaf52Yu7qx1wFMBiQT1iOJeC7KjYzjiRdYuWA
LAHgu3F8aAxMxKsRkUWPBfq/c4wrPCA2nfR8WSDpRnha3Smi+JOiPH+RECY5lIqgca9WGEzTELM4
F4UzxZQePKt8n5TfqUzVlQuyW8DA+2OEcDSxic9rOaT/IOATybs+9NFZS8QMz4GDEhIjA0+fkshy
kKJDNAKMOeb3ofKGh3VaKleYHqs9LW9NvA0EGDx8LXvg507dtQoRbfoZhfnwA2FCk++2clKh7nv4
rDCbX3jIaarJYecPFul6VmZYPYY4i6nSeGviJKSVeYbjMK5jqnntPB05aR7IhQndde7nVRnbDzij
NOwHd4WMJWeoBTgOAcsI8Np/ZTELC3y6vlzPcQlBULsughjIt8CRHETFL/dMG6AIdlhAR1R/3N9d
qEr1ZrPyTINXf/hAGLqyfDIjxgSyR9zVefvn7gZrd2Il/QUACiM5+asxlnACWJdwt9w+lQv/lpek
GaUaDJnm9C/DAWTfXD1QW4L9bOdaERyxRbDeUW90ygF2QoH4IuYuxfzgdJRsk000i8TOQHxg0UdO
9OYiNn/uGzHKRo8fTnFeYkf9fjUMVABBMX3MYG9lG7KHX+fyOAI+HLmy/nMnjdfxxPdnzNUwtCkC
OIyxMBL2J0I+UEek4nmbtOkZWBUyHoNOf3bIc+Bd8hiUGGtKvABmpVgv8IRKRtGJOwD8TJQrdsPC
wpzClHsVOjpBjuWV/Yf8VMv3Ac7L+mlGruN2EwLpvzgqxR+zEYsfoecoe4z767AhmFO4O3UFCSSd
3gEGipGvSkECRjqvfJV07Qvxv38I5WcybODSBmpT0eLQOoTajNn6m9t9SlgmzHZTQXL/VGqiWBm5
HTtg26XDJpa7GIoJnVzYTBO2bwXqE5ZdlkIYgwp4Qjcl+diE3tEomyVYiS1g3pcVudg2kpO1GH6G
ummRnmVqXKgroswCcRsofHHFqTjpEVrEduzWPNq8cpGbTJ40sayxss6Ni8CVHpHfOhYmJcEHm8ub
sNfMYgeG+tku6gHpdC0sl1tRvD/OHpBZHigxQssS8MlQlrhYddylVwkJX8At+mikH3kDZcEeDeZm
23vg1GdJPvu8bDqOQgFb+HUtVHxhjU/8M8oh9bNE7fw2Bnyl34jq365FapLozAcqE6gVfcymm1bE
01whAADODTU/v4ZCnMg4uD8WzdtzTJviI3OmAke9EHtOUmIKAXjb/wgN+iXKg6EvWPc3HMzW28QC
1/DSDjh2gzCMDp1Hs41X4AVwzia1BqVMLUmLtoK4MHpTl9ZnfbPDQO7tC4FcKLHlkiZVWaBTaZvp
cmLZbJjRkH8gfUbQlAIbsCG+YwEdn31k4EUNRtIRR1IXBKgQZs9rNBLuSkY0gcrOLmT+voFlJEtd
n43+CwW8VNCBMGBtUHgaiYEXPz7cyygFeRz2uIszTGr0XDDqB7KmNJaekTVdHArVVceTe9pdBEF7
SFcQazA1ETKry8981g9RkZzA7hXk/DPZ4TUcA+q8uJSI3SkAZp4Y38zsO/Nl8d90pj8g2sSG5zeP
0kyCBldwADqjYPbGi/nrnLQTqOYrH1ufwxRof46OheVL3VXLrwQMFDytDX8qF2FbwtWkAppkr/EO
VaFduk5pnB/66aK/1+SjCjZGea8dYw8+OGUi3pKluaLkzG4LREZMH9NYtPLeLR86Yen81yMQ8yQ7
FkOJso0zK+GOMfq8CPQOp0r7ihNgLMVHLod26H3y3amJLLryN0qjk8wEHLwskkZqFXs2irIk7EcW
FmFJeHNA5ybkylCrai8ajdvUzRZZJGt1tPnWWgRK4c7HEAzFwUzTb0EzbzvC0h70kZoeCa7N0WJq
U5n/QzLAiSg/GHXjmSfufwiHoewrm7gzk/A9AWSBBkDrAPY50XjXo6sXSPec+mY4t/DnsoEC+4pg
On4iaCcGlS6Z+j5XieHNBYKtdGcY88RJG1SPS+1MxKYz9cOTevbsKcjPoKfRg3owgqxn4cxHZMZ3
2yBOOq7zUIyzuNOOzIRiZUUzIQfrVIvDPwyYiZEersAsrjpKT2eazSqMXGjF28qVWtXSmqcL5LyQ
c3O/Sjr5b/CXjs0EsNSaSR809Uhl3HpEAL/9tV08AxNrm8mu0EWpIKUBaJApM3E6kh5p/pwXPvFf
0UuAnB1VwRBCz0wrDlVAdoRbxLyPYD/v1P6FaifM82w0fnEo8Ih3Amllyygq+s5ZqPShQeZhBrfm
L3OnVcyymGsBKIXI+3KQ8gXDue+HRl3sUog0Uh8nl3lijhKGKEOnuth8AwKe5uSNwiSBp7rmUH2m
fvsYCb1O5k8+XEKzoHUAAUsOcvVn+jxOLSLIFWmlF1Ye6wfp0GMAL+qnqAEypRd5nz8Y+spmfBWt
mSBEzX35rykkos09aJ2koKrzXtUc+WuxDIzMS9kIoIp3+Ok53ceRYOxynm5HZH6GI8xty844fMcm
+Jkft1BmReoIXSJfERAGFOKQ5DiHwvEdn7er9ZZBzZiUQC7DDuGMrbCCcZBCH10qWSN768z/aVyO
Rv6LAfsylnITSJD5HOBKTpIX0oKsnJrhA8D1rXzEX6TGbog/ic7bUqg5z9udHFTpspXmjDGvmLo1
A6DTCkHFQgkjegmGwFiptBO52k3MlksPhr3qyTokzatsYqx1Vff9owNbjDfF0A2Ltjf+2TGwNo8T
JnPBr5FGKoWUhEK9QCFXW7Vv3Tt15OTuxKthwb09f+ltMW4gvTBJ0y+KmifNnDWr3j2DKTq7vq7u
GGtq0yeykp+IT+VVxEOAfa8rHzePfMByRoXyOJu92UF4AiQ/qghLTFEFlGxKtzfCly5ssYcv11B8
AH7tw2ec0fOdQ6TLTLcla95MFigTbzMob1AlxWuXpbR1LpMsUlbyIq7daAu/8amL1+O9HEe+qiVd
F1bAo8HwSzhV38Fcr5jx25NcTiMP+9q+qYQu1fmrKXcZ6i2KobjwKSFJfbjePORSbtCeX84l7v5G
Z86ZngIuMURv40kVzq98DQxjCvq9mJV+2yvzm60Nay0Gn2BxyszCZjrQfbuUi24KCVYXpPfhFLBz
7HjyP41/dA/YtuqGmHGYv+VEELp4EtCNFSQg+hUe+4tqD5yl+KOLrnf5or3wJCG80ybfE9oAoMSZ
WU045LjhJja+BSjHuK+GV4DTnMy+p0Ek8JPI9kTTvWb9thMcJDMFGL8S+jtStNbHKFTKuWR05SPI
tub5MbuQmPPUnL8CBzoZXJJg9R9sJj5XK+GdzCO+beNphtC2BwzHUrACRKgRJvq3cQJVSK/LUtpL
hNXedxK7p2Xjx4svKIpCGb3dKQVGgecKyGX9M5CKTUJ8Dm2QOMUaSqd2K/MzVAVuWclaoaILr5dn
FB+LX5x9/YdtYPtpl6hn5MjkpU86xRCx1N/qADuDhYg87lYK8EJoCNb9Td/V3u0KtL3J1DXzboHW
nIToSnUOW6/VwSBOq2PRie9kYWHs6YxJINeWB4lGDOs8N6qitH57Rj/GRiImZCBk8plA8ejfXcPk
NlpAn9O82M+Q2YQuwtLsiR3nqg1dfHkqhg/oLEM9ZvCb3uuGw2SogalOoEWCSaxqX4bvYyhjeGB5
wYA7RrWPgvMDBWcqAPgctKA1E4pb3MQK+lQXHigoAHJythFej1iYZ/IjHBo73LNnXVByHmpqUPie
FFEDFC4dLL8g+VYSyN00Wl4IUfbBxzxlBqsX4L3Fsyf1ZennUcEh0D0h6l0Fez5mqsipzBdcY8my
Vjqu3L89gXOmP15gr6AJsBWnA0p7UV7vQOObB7JroDfis3dbs9AK/HXEMEMBIou7zwwO1w1sfALo
vNyqCwS6VTQMCzzNMhRlDx0Jjd04JUz4Kvt0UppEOHMIrduTmt5pUtf1hK6bFKgP7XlbEC2yzp30
VUBE1UVfzyhs8dXKN9yCDGZ3LzL1oa9YCPuGZLC0DefufB2bcqm0SCQ4rrX3PDl3FMESbHOxNQNp
YJ4oQ4xG/8rD0oWSMKS6XC+2CjUg7Ss73iLDUsEflittCUrQDZtX0L4FB61y41VcCDxEQ0zAKpIO
I8J3IPs3R1BSXz5cM5CmqLgaQAoDAlCCeQb0M8wUkoSwqGzA3lNGAkr4Pp2GRrgfj7TFCSzSaqdJ
NJOHCcujQeVBv5eKZFYigVUp7V57VDT4hNm8kKRCt0sIBslo/AoPyxh6GENQMqBb/8Olim+nIUWA
2tG98hDprwmIZfLNq8ocYkfmVOuFMKVexEeaUv43BzNhRSOMFBgEqkB8LL8abp33hZapMS077Cyo
aQgddzIcoFohjGuhMsEOO75dF56iSpAko6FBH7c2RF9VDNry7Ov+cNw+bl3q4SFzpTfhAp9J62/A
PDaP6aGKHhfhNSE0NPQyGhfQRwPVd5W/xXoYrbC+uH4Hs3K58oLwXw9myHSnsdKBOo+Ca/GEf/4H
TDorTsc/4BaNKtg2MxJbSyxy4ZwS3LNzIoLMrrLVcEcLXSwFuuWACVDCake2MBzhBjogReJYi2Qn
+BYSNQbE3zJpERm5qyBiok5RDY6FiLhbsvqfz0989r7dwif537h+YGv0SC1n6BqzohxH281Nql/s
qcwp0fKT+1b1GKPw78tmV2G4sIxOnWELUo0AbDenIvNgh3DPoX4pu+FhRT6gwsX15UkAdZl38TBS
0d0SCJPRjYgY7rGWdlpoOftW90cdO+t46H8Kq/+Hw+IEeV1ecMGwVNJEz84X/6HZArgx7rv/HmLr
pvB6DKCeCv0wis8YBlM4mN3gnkKWI2+1y5+wGnpjMeUKrBsWS0i0LJsGAdRAMUsqzLgcJHRPV9aO
uY23N25vKAh4q300abW+uATCOuMndYQGLqDCVDKw44KtO3OxHG/ZR4kB8DFbIUMd520Kmrlrl9N9
IGtCpBGv+DFozrF3PY3TK/CagQPQmeIrGxTV/2NcCRXV7oS6zMBjnPh63RrIbeC4NmhAnsN7m0n9
nfn0hHtPT+kXXB3Bv4ZpJ7e8w7R7bnF+cRUHsJmZeONW6BPKvgZO+/opg0PnFP0YcNUCV5FX2NMR
lSPLsB58WiUhYUeE07/fzJnx3ibD3smx81pzsLGaFW86WvOpxdnx7SOtEehuyZlfpXbpiCrLiIZh
F6p6arDtTggWyiQuBRQLjLk7i8T5oPbz9kSSti8qMhzHJuWk+ViO4z+816YNIrwjWbGHfye4nnsr
1BOfrYak9Fnvm9Xl2+TXj3SBWxXBjKq0iuWpP998RZwZ7cydbuDuSox+1xUeYSrx6sXPJnEw7hDf
ViWmvVyZhLRSnpE7CGajyTzj6D4DtRz8asH++9QhOzB4Ym5jZNfcUZridTWPdcI4aAhODyRRNeQg
wokbefcQ3+uMjMZdGvQjUg1+U4x2qwSQ/U8uD/4vQdHIcBEWXrcsGThQ659VtWfctCLGFhoOTX2z
x4v+mQZ3tEbY8FTMsuDFeQxYGAdU5oek8YNF9T9WHYtpIQmSu6SQxrXbFF3HjUNHdOpGBV2jS8+3
UWpDbDP2yGBTxssJPJDt8+z4CaDbNVtNMy4RL5f/kaUbbYBPK93WQLdyzQ6m6c2Mt7cVL3ZE8v8N
3aMTA/WFcOcYl5ktjeRkd+iQfaTo1yXyKYbAyCkprOBJ8CfQZLISx7VRK4cjJyYqvFDHSdbRh8KJ
LIqh78ygqkh1bXBdhOmHJYzMxoqeYeEzxHrjSY9OdcS8WCwrR2cdKLfaIFhRNE84S/6dCva11Tbm
S86ImS8mwRv3DkrwQoM1BPMJEQ0KKkqHIslay8VJX1L6BonQVzOVNrYdlwsOwyBF4P+YGRnTx+TH
IxO+dimGORC+WgimixY401Qbmsc44iPMhjHOxhhnxeM5CiO1vVwwZNwA+xI4+4ey/7v7toQHxEXd
EC2V8gb6riXIs1PMWQJaHdu7/EanQYoFDfKzx47V31eLLrzlCc6wMIiGGJUxJD4lcllBZk8i0xi4
FKA/1mhUmg2zpxgca5qkgTZrXIgAYrt/Lr5JRu9YUI0URQltu14Y32VEPGQ2IdF4tMMH2vOsRCEw
u+HYcqtMLpew3mcoQ+oILb0a7kaUGSxvol2KNQhhJFR3mjSV88gaYG6psatRBY1IdsGU/wI5z1Vu
sSThfdhEQVyruFBT/5eKaS/yYY6Y8Tl9sy9coYPrOXlC8iLKup6YIPhOrUMjE7jL1J+BBCL9R9IM
PVFtzT9Hz4xapHIhNYsQ38bLW3FB2EmfIBGVn2CSGH6/f1lYvk3Ijy+pANkqvOlSD3ZINKxnFm7k
Rr3W8xsj6l768uWQwluIoRmruV6c9Vj1nyxWi369AoyWoK1J82UYgVBQdKjIu0M9wGKEkuEOaVNU
fLWLXTdlqU7zBS0G1rQhjyNq4YuiZIkjyPPW31OWeehdfOMFkIzJ/s+m8WyfFctB6gIJisXWdhio
PHhh7m23Qwu+Qx9xjux1iiQ4+vS6wDhIiMn6ALKgkRD9ycPdQTJrXI7+9VBtKJzUVGSzodsgmS7s
d6JgWG+/V+Vvo4ark1/b3FnyjsQNuTd+NB70aIQqsELkkEGhKzouwXaNGEv/1bfdI9DfND6+yQnB
A6hVbc1+BrvlVap5Ku6cAlp2PRkOgXXkaXJ9/kwcyUHTWalsxWg7Oanb62cv5Htb9YuXcToiWaJt
2QrTzIqhW8oXZ7r/PBLaAE6TLY35OaYFNsEgD6Q/bGADnD9PrAHGxRI6wJWOCBI4RE+sL/SfTYM1
n9kHT0cgDtBH9Xs3AetsCdQTdopbTOde+kBMSO8Bm/c7aPbAalOj9Y5sf3aYqnfVsr14gO4YZ0hz
OmhS1mgGSvR+5vNM3A6V2CXi8FEKZ/hcPS+2hQUt3aJ4QxeHZivZpT1uvX3Ux4QKNCZiz6ZXfCLS
ec1K5InDIjp9WccwucqdOd6efvL/OJerLqf5BmrgWfgrwDqkukZV7qXC98QqCJTHjpErumurLCjE
5oDoqZTeaLDw5htdvVp8wO8TeFkBKCHZdoY7GA1TLS7N4O/QaSmU80G2JpoQu3Ntxu6BQMvGKbae
zLIMALLGdtQIb5/pdk63Yjr3O9rgA4hGaQcIpixqepkP56IG+J+TvW1a0m63Gqxu+1G1h+9ndfU+
7JmZH7Zjbte4lM8UDuvQPYcnr9ku2AmHsKZOPe9Ku5J3/mUy6qa8cBwogE1Mtfyay/PBRwJzo5D2
Uq+RJ3nUk9NY8qguMib1HHZfe7TbFPRW6Vt5wm6aYUn+5skuJjU+8seXiEETQtQxFqx0MsX5cNnP
+QWALNSGDUXnAv5xpDCDWEdJEc1LpXpyiw0gE35HJegBYN68SmQXHe6qZnX+UgTBUq8EU0eyBXb/
aRpjRDIcjJCCwpQ55lIyZmjvpfXWc8+LXoHWIBrKVayIgu1M7QYq/MxrJDV+rzXJQpC29K48CM6b
MNZWzgjxekKBH3POopXHDZLFBGggDY/Y6dND7gLbdkhq1l5f3B4s8vmgi9Y+GMIljMUU0kZfEt0x
T7q8rRyKeIKKgDCn8NjURCR2I/NL9tNiwPWMSTglan9chCm7jMrQVrYlomT8sRm8L2ewPXGHaAC8
/T/jdheEKbpjzWs4HGjxGXI6x54kYK/uHrQqJrEx7JI0FggiBKs2VwcvgQFgLdQ+InYJEXV4Z5WA
LEU9UjwYJgvO6/Jm7T6qNvHSq34S3D0rZByewbvnoNPKM0ctKIVnpWt7TZO8NtIHgf0DLvzy7vQY
bupqdzAJC7AuTidexCP90UxkawRJA3ebGZHROMDfSqaMO5BnzFmiJvs2+PRw5F+0Ly2A5i4JJOoq
cGNpVJ0gNiEvRLtXN/SBltNz8HcQP2vmyY2x0fFEybBdm1+TtaMAHNsxXQjp8I41xuoE6Apj7tDW
Z4EXOJjwa5PqakPsATC/8otQ9DkvVMHgb0fCCl9yljqqfiMz79FeTEXvswtW4HRD5hjOUjRWy9z1
UHEt5NexXUgalvjipKUuwmMPitYvdcvi/vFuPB+LuMnQmhfXiGLAgQi2Qhf3uzOFCsQ82SsyA/zl
bl3yQ3+dlqBvO5nf1BhoTCu0BdYtS4K8/EWBuc36BL2rRKYtjJRnzK+LwvVq93MpIiLROHn9/vlR
AZq4vtYYZR49EzebFHB3i5Iu5GgEUFGFRQGTHQK1IGPfbPz6KgDm20CArKwqMhaxRhsbNFOGuOtt
WWsC4jmnP10FjWdVSqBaJFz4wFcAsL5Zp1poAxpPPNAoqmwagU/PNoUfSI/0wurK3jW0CzSnqp8z
JUIb57ITGdcSyXu4UiO9rBMVo7bmyknZIr/AzUzwYjzNUztNWuWN3QrQ3SIMMBucDrbtXzd/cy84
uhFtolY6e5lyBq2h83Dt/5A8kNG/36kBc2KoLjdxO2UiB2N7+MPjhx5M/C/Yhk+eVMKGqxnZbeP0
aZv0RuawpeHID40s7hPW4z3YJ0laJVf62+NTmYjYb+aPKDptNzkQBtazaZfzY9P71qsoh/PPwugT
VOQLkHHJa5OkQTP0+7G97wUw55GnNTEkErIOP62cZj9Z6oAUVVc3r+hzkbJBRY8pyKBh0fVIMD8G
b8n1mWnmePdBlSv/aj8x5UXZW1Y/mlRNVL0BPTweZOQTOCoSpAQ0/sjGuM4Eicgmeb2qTB+YudSv
bWsC8h9Iakz9ZmgZpkdGW/iEv/3kUq/lPcBXaz1kFoX5FKWY+FrJIZmqBjpCrotgcXjQmxATjZTS
OJrSJ1h3qFEEzHAJfSNE24zlD0lHP39v/1MAI+ahDxMydLQ3FIqgI8NqlaNr6bYCBSV90vWazarZ
1wY47n5G/771VyNXr6VlGAjqRQjv2fnLO7dysar9IoRKqwBuSZ8tnsOhIUS3HGo8H35laZClo/Y/
8OgDNMP5Uj865RnU8jbFraGQ/Ppni0W0HS9xe9G99LtHclgIDy72LHAw9YSe3DB22cHrudxATLrX
N5XA3VyenuZpUJRb2M/yK4GYZkKWfZAmwZJsZbaD6452VhsduQoDnwOnDruGT4emWGI/uzQcKrmJ
PrHfziP+r4xsMPPx5c2Lo3lYi5FJPSterb3FIYF0Ujfom00vBUIYvHkHfN8CEN++V2Ih3TMlF3Zq
wFDUjjNqyPGKB+frgSJbImb06SPNjJ1yDniJmLgShQGNpFqtKIMyF8pGa1gNJ1Z+WFR++YcVSapr
BFFfFgsTF3FSOVpc2p2Z2PKn39BsscP9riboDjSUYStPlBaK0Wjq9vNttM+fyjf2YM+f5mzo8QT5
/k0qSK1lArBlBxxvNQ4h2YJm3qtn3hvsrlFCXn+FSPunAeQzJI7JLIiCalPPCmScmZLy9aI+7su1
WNw0W1Mt2Qf9rfjsKaOEy0VrKp/rZX3S95qYfA6SusjZeqzEfMp3by8f1bDpt7gEWohHLlOGWbXz
g8ugwXiQKjuh8BXjQeRDuHC+Iod//O4NcKOZS5npmQAe2gg06aOPyXf56rUyx0YQncDeN0gq/nZp
aeYNwZIGgCQrg5sBT6Gm26e8guWXyfn6ABsQXl7TNl2lhBT8kEMnPEp/LLqZMM/6Sx3dYxektuoM
ZawHOJoohIQ5BINRNddU/7eLbzRM0rvWF/gbva9MRWnsaoJBkclSSWN+KA0wqkAQPdmHatj0USzo
FC/ZqDCMt8dpGv5VIraoAUwXJkU3dX5NCJMGYpUGYY152v4TOlngKHtKUpjXGi11d7MJrwH4UzMh
b/sV1t6RncDg8O1X4eqiebmhvPmR5VCdcsP1BzK/nM80gDzzp0WMdIqd3HrgMyDuV6TbpZZq5LtQ
n/L4baUsKM3TPsrUoH1Zbvuijs17K9BMFWS8MjZsN6A6kCu0SG/eqU02FkbO175OfgZoF4KRvMAw
QMexlFDKpH5pqJduW7uPmLESfdCovCcjZFI9NV+71/QdnanbfnJaVqZHVSzlIDywS+Qlz1TFpqLC
/MnBG97ktrnjZcQEY4Cz4TvTrs8NPUVUus0C50hvu02O6JaxbnQcylsjkUYWJvdGGQg2ei5VLZyZ
EpOwjQcBSVZwk2b/ihfFqyMhvmkwvaQ3Ma+Hdk/TwzU4BbEsMkx3OoflvV837rXarW0+uyyUsFAB
fvUs+moFuWVNui4YfLKrVSuQluRbsbNBFtFYHSIKjoN5A6AaN0gc7Cikeud8ivfdmfgdqR+bGeHz
RsdUR8C79/GACMAZKsmmUSIbTbawELdxem4e6Fajy+CYqdtcC/lMwPG5yOEZnZ0nF500KROPN1VU
Ka6UC4fOdsq0PEsFe9k0SgX7iGQzQJHge6Ig926l7n/nOtKT+KhnOVbV7Ww1T/XXBcFBeM3whzUG
qzLiORoxmmdT18K9VOK/pwhbBukIDpNT9TRMsVTUjCiLaGALlKA/kiPmAHSub5vrS1tEQ7rmg8q6
R+KzvVHBB+97OQP7axOMCQvQTix2E3vFbOvuWaL3mzxEeslhK1XK6oZq3vzdIzna+cVyb/bO5XBu
IQwxNy9NtdoyPP7qIe000MATn3suFl6Xe17gflrE9PLhTveNGb3YfPff0BJo2X3rR0CRea1duKlq
9UhW0hi4GmVLMIwpByXMPuPnjmqJOil+29qDvqjtFX4V92YF3qSOU5ap8p+vxLdze45PaFr/2J/e
U/zZ5Q+nqSg8l1CGZUgkUDLoVDrVCiZu1pHqSmRePwUPAkxCha/KSiCqIQf2oKPvaC2Ygkr0qpXe
5XeD3adQSmtBzpP2EM0O4+s6PYyx7SC9t98Gi/hCXSkYwLQAaMUWUJG/MEirNm44NrenFTct226e
xzU1o5BUUpQVXVJbRuZ/5GWhb9cqOqnsZDon8lpzy2YHagLlcIUQUknikNP3d7YvAIHOMf8IS+q0
PHp6pmmSvynJWGBIS0UB7Yc7WNI90eF3P1fGHKJYyH2ip/TMZOGwgLvO0eGqobin+6S/WWCAYtFR
YpVUT9PD/9DXFI0xt1SKRxl37669tXemYzrzt2KO8PO7jQSG+jDg6XftBvPBF9Le8tLCORsHgPhv
YRoneyIHmOfzHBVOzlNh9I1dpzFLyAWixT90hDNFWHuhCRdaDVaGsxoOlhW+XDcvCuzwraLEttOs
8RfGyIaOYeUrtgj/sM3ZPd5kaJ+8AA4VgBtAqDG8FQk0Zud2FA/AXEmKOoUgiNIkzmSxKCpNZTM1
9NMMG/ElvZrcihtxB55YAyP5a0Fcmbz9NOvpka9KfRR2dugP9fUzAn7JXAr+gJkcbh3Utj8ZjpOu
FLZeY+Qv8qBAlqQIXh0IOzQwfbLB2gyaBWFtq9SZHbUjrmHR2wNgjpSeOi90FFgnOrvaJJdlkXnC
aasj8PU11/P6Yw8+rnTzp5Pxu3kTkG2YLoJsu5QCJelpbrrtzhI+ZHd7Erabl7t77DhaqRJ4IecS
sTfvmNO9jsNirIk4GLtiSb5Rl4ojmxa3c8gxZX4jzvhCfpXOPSffLARY0CTWEfarV62BHgqkcYyX
iPWBopX57iR5x6oAu7Sz5LyClwvZxkYc0jpaczKPzbUqhGkeOLiavQj8hJlzX72z7XggyqcEODjL
sRdhfUwnbSxULSo6F3vs7J354crMnnddBN8RK+r8lnYfC7HVE5xFot7203FPq/wiJh4sSdhvCQVq
Jectd0R1yG6bPduZhAZJR0WPxHyzifuitJ0h8a9tWFnD0qZWT1tuNefxFBf5nfA8zq4z/iz1l0ZO
d9Q2FPa82/hSIYbAIeEslLt4C+MdFG1Yd52ZCPoTy1DgGOJfEEasjEx80BId7iAXXYXVv5uJIRuh
j/E0a3K/Mn27JaW236rM4wpeEr1YC4858A/5GuskkWb5yGq7vlzvUOQLu80ZTKyhcCWD38T54ONc
SNnDoUb3gUWG13aGyYF1ILNqvRg3TWCV5ku1R083oau1FIcaoTiqA215C2zhT/a8FO4ydaJOdWwC
fvETOG/kj1Z7/nEYs2G18k6JmkFHR4+zwVqJu0DR974wNDjk/o8lOU/OZuASJVxAU28vry8o22GI
Rtm8FzCRDy530dghsRRvqldVugxeVGTPEmETQXPqS6epb3ciltdQkjMyzYcs3wcVocCYZm69Kvdu
0dLg/Ye+bsR5EM5bQY4N5ySxSVymQBHjRDJ/Rx1f4tKBCLfYySslEIlBKm4P7x2uKBhGOIDwFivR
DZCEGtWrkJ8vfcVz0EOuPT7ARzyaiEoOYau2EkFxmyP9V+iWc3zWI1RzXf/KwtluO2GZDTLXFIYv
a0+qA2/FjAFYtkkmkk1w6uiVR3kcWXnIfoQc9bs+SIJzx6q3Mf7sb3sZNIY2UJZtXGPjQjnCT8eh
ChHi4ZW5mh/vLwmWZ/EdIeFvSjiVmXyJWuApWl30N3I4yp0R4JrjrYn30I+BzwIo2TSkbqev34aP
vRKWyVWJ7sCSqjOeFcFELQGY/8jkfCWCwsPHifZpmn5ERdrBzlpD9QZrSyWXw3xmshKIcx1ft/r+
7M2efcge+qLIPwoIchLvCYMQDPiXtJTIuaH8vCNvejw7e2+4V/+/wYglYBjcJsUuxwqIhFPyV08e
GezkieHtIgCGO3ItpMj9mq1Lc015RN2+rhMeEKwdcXYCUheN6NQHMYbF15jUtUlPXPoJ6K0B6+vX
PFciPOaciTuNymcc4ebn22vZJvG88JK82NCk9sFnZ41O+vg6mwzKjD67wi4iYtJXgbXDf+4iNPS5
aMigX6yOFw8By9lC3g6U2UqlQUU+qzmdNZcs126xMoG8S17QG/ENkRFqiQJJY7NLmQl0E7x7Ld6Y
qdsWM/Sdlihiw5hjAkxNTt3Y4c5LoRUOT+cdzIKSEs7FRLjKorckQrlTSczk8OXBWd0hAgvBdzOQ
1MFO1oNvlZm4S/BjwoJ1Jrx9kDwWdRth8gvqGwzwaeDWcM0vs6SL1NhTdBTSFYuv00701qmbVUE+
VODo0tGuutqnPbB39HwywH2aZlHKP5grzvrCd3/BXOSEVHHDjXPDXx7HZfNTNyk0d8EwvVuNmdHh
0i2cT6bjr8/vxSv7C+nIjx22ILor0nBpvbfwUH63VZe+B+5yaVylqT9T+EQgkYJ/tcvwpfAqC5n8
cyqlrwgDKkoIjwNgGQrcKRz4DyG+HLByZqxpzvkr1HDwot4NVFCSJAIQJkH3xsNoo7Y5hQ1ap8xf
Py+sRO50NZfc/pEbLaMjPdERK6Vpn4EWMqHTUCHm/mHqbQKtkzlBsEIJcc9Z0riMsPOGTuj0vsKE
/z3xUUyU8WLewbiqzFYrPhUJDwJ0kXABzuTWP4PFl1TGSuVM/HFTreeR5kIdx0VDsm2Z21EI0PDJ
bwy5veG2JIpDCIDdWLy5BYSIxq3TUfg+83yHMZQ1cqAgTGT1oLqoDkEbHtujTSuzssyKtJfRHAv4
Da3VeEhl+VmVyVq1gyDjsZzWSZOLo3pW2OG7YQK8+YM+t+FGTimZEFexCecaDjDzPFK4dgZhqVUd
goyX/e1UzoX5r+C+GStgXlnrlfiinBMz3wkafukP37AbI3drz5zSsXyY2bdEIdKgmP0NmIVHIxdT
MvPLaMBDFuYOxpE7yCyqOywNyLFTC7V6sOziwoT91mB97IAzPP3l8KNSTWHUxevqgvVV/j2y5BuA
1/XRsMjOxukiTD6EpudEpe/2HIHyDi4MPrhWWo3LG9TfTrkl4/RV00mwCGqeke0APa1k4ObI37x2
13X94b42eupr3LqKg1TbbNQA4WuCVrssKAfV0/sBO13ZItne1E+1DQhwjnahT4bGT1T9bxLST1wR
LiBae/lFqPnWjpghBnoG5cx99nMw18XV+MIU61RG4LNSvAvNlUy+xOnJo9SbBz2GwrWziq6JxNzT
B/tIyy88fa0KyUU0BxhkYz/PRokLD2Un2TxpRazslFAVwJ56UPh0EhPq/tQ5wKcOXma0QLoLc7PX
0uRPtxBFGlNx/2mirQPUuIMcVGL9jO+FAAD7iS2RUrTfuIR+crXJhUOOytf2rS0ef1FMrIFGbtWd
wyknbU+LcMJdjKby5tdU2EcsJacZgwGiQjhd5Rxlt+JIexROf/4qQvA4T0Axc3EgdYkJXMjCt1ff
QySugWDHB2WhxsowthEH3kyc4fF00BfyOqyYR7LIMviUrpEaPydgKPSp8r2gyi4eb/Xsix2tARJr
S3z88SAqJ6LmzocgoIc5j8RnfIST1BiP4OuZL6pbIoZt3RF8y7aHCqAkAeD8mugrrnQAO/B5AQz4
kWNzajY8mXTU1bBNRmbPbnHsS8A892CQSc8itQ3ChbMvEjo47SZsj7P4siPCFU2sW59jz+ktiXFn
ZljS6HH2JCPirhIlu3rjsDm3/T0rESEMykZO+My+LBGwu7GS2m+9y1Rp4iBYBnBxfC9JxnaviGuu
CSFL3dB5goREJtLWtmUePUHykHVoZUSwANoae+zWI5DV3GDtM5HA669TR+ad4k0mmUDnBuZoCYOH
fXGB+ZareGqYgfxNHCBuFDxJ9O/kcYvDJo4RxiTVXiEN0KtZI1G2nTHR7xXQ3DQswD5neqSXeoTf
V+u/r3dKlv2WPCcOJzi5ITS8jpaUdoUrpgBQtyRgnV6LxYJW3yReqLUC8ZCyg1ZzfYZQJDxOL9lk
yy9URvOzNPxnE4zwrgPnaxYcF0gikJBRU8lBTfZnBJM7Eg4D5yXCO+XqYrDXaE5jeIfwKC+hfnvO
AAlkDq98HB1z69mYYrlIZeuZ1LBS4CZFcefsJ7Ambj2szz5ky4C7ENuCmDg5p8MAS9rva9DShuAQ
6KBensviZasuUJtwAMgleueRbL5KvrOZH46Ybtg4QSEOrVXNR5x88W1njcbn6bRukv810CmpUHHB
E6Vz+R9xUDwmryViX+L67z4Ie/UdtxtvKkvNJU+i/USvIaJ6pn+sEK9felL3Mx3IyjzKkz5vT3Is
zK8ZZJ4goIARu5Ww8eL4w8RI91hZJv7zv9S1lyur6Gzbre2al+GW6ZkHIKb6OyR7fdjOysLb2LVb
qh5IiiXL/k9X/t6E0U11rfx/KPxGB7FE9LiafKMKmDNbG/ggIz36/0DED/3hO7spsQI3wSEiCIHR
cQs6CsUyk00fzGoTI8+2ftV2VjbfxhO4bfYuQzbvKX7++wG8hzUm79dteQJoEDnErpzDFngVJTLu
9iiMQc7OpT4OiOvxQunrBc1lTBJFJ05NQvbfWCCHIbMqvapVIkeOiZ9Et3FukctSUqirlg9BpMbl
UiGnOQJc+kNF9za2CkqjCQ28C1O7TXg+dYUbzJWDEu5KvJInBAB2DXpsjqn9Fvyt+23oGE5R821g
X9FV8fdTLIKaJL5GplTo4Nj8RIqy9i5xQoJsmQlvipnkdkC4cRB+5hRuiEiueKh1QyAfERwQAwRB
u0yncyaw4hVmroDBvad/rfeWPUjsqU/k5A0AUUR3HNJNpi6fayZ+R095ArgGno4HOBnTqQT2DAB3
Fw7b27KQvIRMcGAHtobs/KpbSaBnn9wW8wMJhqukZbyDBBZKnhTj2zRAJNVuyINgXpCkenYJWM0W
hryymJHpJvdMln5VovptxFefI+RtVWZwsj/pb55UA0DPCEnYG/5HoLeceyAP179ssrLfowsrBCZn
emg07wk7iRNVPb9xb9GQnrS4ob4/G4Ye1feXSR/9bhmjFaPRlHgPSTN/sSNR+rLyyVWSj6YSu9X7
randF97mmr7M3TxhBLvzu91WSy5V+I+cvg4mG/3L9myDphYWWp2elE4Q27ByhZ0XGsc6CTUA5ml5
tHvwXIvY0XWr+NpuyY/+KERQVzcTLZd4G72DqgNGHdRNoP0BSl3MXYxIZP0KuBAiCyptDjHHZi0x
EkhKs3DqcQl7T4w73IUpZqweVDpYafvq9VpdVsvbxOoEefcdoVKyyNkJko5r6/C/OO/QGcNuWDpu
FQUo57IJB6N6uYHrT4w2/4gtGWxjPQXD7WOzNFQanpUs0bF+Wa6sIh7MbMZt4hnHum69DcpHj2Ky
tGwwnO8/wnILAir74jzlPaJewZP+Ahn/pHgO0myl9EdWhHZ3+zFBMUjcJSAD3pt2aLfUhqXbytNg
FcY3cSoANxVQPs+PAi4R0pcg5kGKBe6faPVLe8EMUPzO2XZqDK8anChB0JS+3hb2H54ZoNqPbpu/
/NdJ8I3u7GEBuyKd1A6KOyhsU7ujsa/SFXR0plJE5DduFRzsCDze49pVaMSArEEcfan4PM3sSFxq
fbwwRDm1MmbOI5c/6Eem0Ul+mOy/xaQ5MXb+vjeCfsvpTScSu5khcgLO2l/MKNYyrMSh1ky27Uts
BH2aCRysf6uZzWa6onmvzVrqW9DvQK4g2SdmOVKJuNf9v6SB1w4EJ/ucwSASanf/XL4rEMCfyvRi
kWojSw/SHLaM1J1Uj8i4jdAY82E9hTqtyDcjR7utItLFa7mq31XlrQ1ZDjdXtCVpVB3/yqUy0m8n
GblZfCaKnaSKOC03rYuNJlgtF2iHZqc//LIB5Iqh6gQkuABY02GS/oYJTzchhB2U8OKmSY5ybdv+
ftycNW1MiPLq7p66F6XaMn7VcwKJ0bzWpTQWNdzNv4q12PtONRJfUVmYCw4yfASK4pNLx6XMeGD2
Ul/ZWoKkCSIYMp3pNZuFQEMou3bX4kRDLPwYr76d49hZmkCg6WO1XWNJZ+ENrq3Nm8YZXp48fpW4
nCIq/WIVNDrM33dFwhy+Dxuzm7FvTQf9AKbxTJcVyFPa8BZ9qBURya6+PS8JFgWrYxT417/YeK5W
sj17zvAoJXx/O/j404eJjpJnBSK2rezTy4hOeK+A4C1zkK1C192IwodaW+qH30Bx40qlPsv7LEfE
pHbvKu4C6NapqYSspx8ch7+RyxnUbrYR3AneB3swnM934Nx1Kh30zSLVtVvJsIDBWkVQv28YeuM7
4qv8qZy7GdPFZoAsbrbX1m98q5l/8THMTL4jaa+B2EmLKepGPR2jfwVPpagFakeSXPoE57zw3oHh
WHpk/LUPrPgHuaV0E1Q87PtL2PLg5ROhU8FeeDMF8wQZwkvtklklTKKdmqhqAsym2SLgH+tIb/py
i0ISupXT6fsl52Zh5YehyDDOPVMTim2MNIjOhruKch3ft4i7td2IS6X/ED038Px6J7AOx4mNLWlY
Xa96SpGznEZBIbyDPfzOLFT8iZFnnsl0r3vcCLFKMWJ9QADIiD/rg6nTk6wuNmQALBW8iTLfjl8O
6rNjjkavoaY5hJwy1SKuvcSC9Ci3linIXyr1TrmdbAoWkzsdNMJcAZvZymDHOyKSO7bdhtMDZiZz
hAgF23MP9utZO0ysekhE/qYkRv1FSuwKQFL+BQLzMQ8NYHLZOO+cXyv37ikhriooTPJa4NMdnMsF
R/niqHEL50fYzy5M9O/ZEWWQhh4QH4bpvrTE1IDgQUXTSZ39AcGUJsK7n748TuPCQ7zPVTklLlxI
wbNGVvtlY1t1hejz+2dQMccS/XAAbDMBcLbarSXaTJ2+WQHmxykiLcxSuQQdX+erWugoKwc5pLYP
oS8YbGbHuEW8VNVFZzYYky9IzwnXHsMm7dhMuBTy09VnoMF1EgjzxHuvdxobuYaWppZRpLIss6FU
E0NNQoybL9I/8JT6b69/JwSEyxsdTVsRUQba0zUzkTepjIjZlFP2+0O2WzE4AX6N5+llsXGPMi2r
f1LbUBt4DgmE/+36czafZweAWEGtdQw+9vaYoACaFP7mWWlGCAExddrOQnpsjSFqoJiyLBPddGeu
XRdzUKj7mVNT6PpNYazwINVzAhvzCcvkR+5CkGsUDbS1MY/x2xeu255QQ4oOcXViSn65UDbPlWh1
tWfVE9bv1DZYmWI5+3TKTA5hD2CEDfJvc9Gb8jvWDn5TKPdWPH8ShBoG05TSEyNxoOzZHdm4F3KN
lheV/2WbEs7sjv5dU8dF24966Xww59g1Xc9Xy65sWEnd7jLvlt/JAO7kOLZLOjOtGEy4lzPxV2Go
zdV3oopxGjDvR5Ano7QasfseiBrv3joarrlENH/3jLgPHJ38MbOdCR8j/L9EAIDCxQDCDbtIaW0q
fwTI1TgK6qc4AGtXhsi6zyxi7IdaXJ4SeM6yI5147QwRNK6AsoJE/zJU8fltuIXyLOtBBnMoyLal
cWIk7gc+Xu5NvnwMkVSxGCaXRhopHuO0cJoMfcafTzgHFCMUb1C+7GFf2buk7tdDqfDnY5iWZmWA
evwg4aRxIMLoxZMjDmFxsPJRcTIsbSaFdv3yK8J8KegV3Wv0nH0GftRqOlO8MrvGnLka52TuD4Bh
ob0A4MDgq9uHKe532nLb4znu8jtR7tyyU40X6imQ8fTBtfxMPA8X8a1wZTSNSwG+ENm15S9EcjOq
CJbkTSEBhNSXyQDd0fVp6Bn16JFdc7RPNXEefwVZwIFnzlwD8W43Xh1pEaEjgQVdb1gnodOMEaCT
7/KVCls7QkyX234QzCPzkTJKzsx6+DjYRZOPIUO8cqVNOKNbJGgG8aDjkj+Etzo6+YeFHSPYJHWY
oydYepgrM+IxjaJvRUV2I85RCKbU/djfc3K7SDBARsWRKs57/gG/pp8qVoyBSxjodl2E9SWy8scd
zpWl9oOkp0k6GGPzhnJyI8uxH1h5ICc06EdnisevqHxdzgmB/b+lmCHqkjjS6G/pGEFVE9Yq+JVZ
KXfhJnwsRSlUvgo62IC++tVYzPfjOuE5e9WrKfFv4HeIM/G6xu2EusR21BocCpgD/5UUBQ5bMppX
lvy+hgW22SHfPPjzwVpA9v7ii5zeSSjQYJyMTCj/qlENoH7jrLHpDPC4BI4Qz00A+H/Y6fl8qqls
Ba//m+fRE3i/RU/1y/dWuEUC/BNv+dLoksIrHInu/HtlyJXOyqBdhss5w0NOSlp7jQWeX+ZQEpMh
rVK2dnldFwxMhxmgrVv3+GGfdGZ0iVSWqHYcXJtNyWPMShkcQFNIYsShJvWWcSNLTezk51Q0RnbQ
yAkecWN6fuNTecntLBCO4ikmc5991u8uhkQSv52bO1yXxQoT8R8sCMTjFpyIm6QaCCJK7Qb97Jb/
BlogD2viqvgQXeXnEoi4qro5XqKXmoNDja6CWMrVJsea+ZwDPP8IOQwoY1q0BZHfXRwENP0ZcZX4
rDSwaXRlnD5eu8P4j5e3/Oo9ycXolC7QgugKmACIVTPgW5Gb6ody9acwiStGdk2Usmrg7xmSjqkp
PxHDmBR9ZsoaB/rtM3jyET7OQfBK3T8GmkU+qFPn7NpuKgu+EpgK/qbp89jnjGrF6AcahxSCYqYu
cvimV2KjSjppGW3SENAKt1hDALJ9q/crILJ4AMJ6WNLXJWkVrkFhVY0vQzAviKpdLqNPIgcNWMu+
c4FHAB2KUEdP63z1iGHM4sDVmZ/P+/PrWCe+Nds7Majh0NphoAyekFq3gVMgvNheqoffOEIfzXIX
ZFiTJ6S/iJuWrqFL3SXPJPBflUS4kvT8U/Zd10VTZ2yT5Y+OW3bDEQSa4UkFxz81IOT6UvyagmGM
ajUtd3a4YTzcJQYUR5DtQhJqszOWIuupHFAAxyU8Ix3y5jXQ1OeFw1l26mkf61+IrukbwIv6I2p3
6+mT4v5ZKF5yqeAnVAY+1VMMZzyV7nwEw63CB6xRDbAKIamXrbw9vlpqY42j9LWBs3rhheT3V+uq
e2NH15l6NUux9OM/1CW14Cumo9Y5JGizgAUS8/On3v8i0exfTevcfHWHZRWetJhQY6c8rEF8x1ZS
MnI1WK7rrhHXYcHkMf+dYiUdgx8sabgG/y0TH2u1Gu4bOX9rB3ECYxIh+F5qh/xeFHzXWxZsGteh
9J0dkaKXIqmSvxheCZx02iUbW49VbKO2Ik4C+zQRTQq2ymZ30HrIGoy0jNHWMw1bNpMRInHX71tw
FiQCELSbt1qOv4uf8QhQk+Q/HZC7Kog9+z/iGEaGojWLdl6BIG78m8ijS5bnGcu6y/ZLAADoB/eL
IvCeed26uZbXkW8GBTng168qco38QRe/QAcdZuTNWfsEWeuygiy8rDASUmlp1i2cgLg4fK6WC5Kz
BkLtjztGBrIP2xmsUf+n0pISKbQ05nT+r9TDOn0qyhzsvise+vlbj9evRnbSNRltorED/afLkYFM
uaw8aJcbqQmw5cQSJAmfOoaSc+eqC9z4ObgSgL1jetHuLPQp7xXOJcPHWpbGGWf4BLtPfTm5W348
d2x0gEvKaVJ5pcj2lMNFuPDdMalPj+Ipf8Gak+5NyqOokwtf/jb5Op0ddlvy7zp9VslD8cJK49TA
TEi9YlI1bOCF28RRzqsIAgeqEfuldhKdIC3bsBnawFcy9yUWOx5ZztSigK1gkiNrgCiyKiqbfxob
hZMitU71djZAOsg81sLk7ultiuZN9yl8BJfGy7TQwTlKpKGGWGLGA6LMlGWGk2xODJGIXA0iIq5P
wY8s/UH+Ub3axekCw0eXwF6mZpVLpn49mDwcPSODWwSabjKEO08ejhUDxeo7uq6p96e49UkAv4dH
fJjvechlj67O4J+YzIzmvMpPwCInuea803FKwVXMjwB1cUaevMK0plM+y2z52dna6O8k++rvo4XC
n9k0IuH95w5SAAqa/56mhi/5WWW294Od0dFsz2mda0Hwc8Fh6n3A6eHGSLmJ16ivo9vNCgPA4zuU
ErXUo3/R8CBuGUD0ie+t4FTVSwQ7DWoF26IhNkhR9vqyNUIEuT+m0clmgokOFrb9Y7UeTWBUj4MG
qq3PyJJWodrrPXr4H9N03IIFgKH5vpfG4uos8/eu+nBNX1wphuADhAwj9aPQkiPFXpV94H9TLWfX
LrVrxSegiyFvtqGNAFuSahX1W83RAjJ9PGOLAUR9BzOebeyDQRJOE95ERY3UpSVisH1dmfrlqHUh
pS5/MOrApyl5PqB81ymrdSQZHaac8/yymuG+3VNvfAqxK1Nl69mCc7xg02dfzTNY6NGVf03QLaqp
K0v6/Q4VVMWzV5buCumtsd1AnY/lMLe7Ela/cuQSFeBWEhCzj7SzvZExH7m/loGHXRiC7ACi/HQu
4H++HUBl3XOq6c3gXdIDxyh3+eXY3m14RcE4B2Int0VbVQ11R4OX4d6Ux2jJhfnqXyHl7k4757A0
r9mMNNvwFwosahiY4lptfqrFb5xS9nAXANZel8/3q/sKqEx/Vk5whitFxF5f0q77kFrLy9pPMbOJ
DXoa/lcCGaNBUuqhlDGQF6+03WZB02lNwGIoKHdYLuIYrFYQLnUTuSfeQBLNmh2Chk9LyjbHIZrT
JF/lOicU+LyU6779eHtqwyvOimcQTDgzqeJkPBj0LIvwI+l6dijGxO64QYE112ZwP3jtvBZTtIhG
+uEsm2P73imNunujeXeti2VXthqjNuyy/SzdIvFoLIbTK5CCkgsDGITSoYuzPfQXmCVyXxBHByYS
Gxxuf6fL/2uWHhmSy1uLwDHcLVXwLfnpl6u3f6iy71uR6k7+JsWHP+zqdrx4EvibcF/jMHyMkh2g
93EfGviMdwT+W7PIdTsvcDBIkP4cnYqPc7S6e+e/uAmc7jFlOego/MZ6Ou2JB+DMv5DL4TChAqca
rBSDtasZce3U4U2hlX+8hCW3mlae8LG/LISlty568rTSSVzziyeqChzjxixzCL4wFEEJHo3rxjUH
ZJgD4xWEn35RrB4mIPDHBEhrlHCvpR0/TWcesqThY47gGMENrc981r/J3LExKE/4sBjYOXlnj1aM
Y9zsX9Y+XDJgU9bk8OjxStIh1wagZO91OXWn0TH6PkadlOWvAtPxgLx4xw3mD76koLw+woE3PrnV
B1IDQaOpLoLbGAe0N1/+bX2FWPhe1/0djuOxXs+rdMdIcOjdh6Seb0z4I5ep9EVCfD+9sIJmT0hg
iSM9lbierNEOxqvFSxITvolWOZ9ODMNX0OpZj4kdT2MLkmDTSdO7EL8TfmzKI9NAUPlg1C6Vuygm
u9t3NvsMHiufFGxdKlSVJyiaE8/frQSIQICJqsPNunOoGeXeIC+utZdNoWyg2nIPo59mU+mZxqlK
qa6Epqe39Tjq/Pq9CkcHUjlZHytd+OKryT8pDfIRzP53E9Guchq3QEInJSqdkuo+npQDGiypQaB+
l4R6T0ncbgl1qqsawhKoB6BSO7F91WtJYb1yd1UiM+tUvBIR4dpsMHJMqHYYF7oX0Ms3Pb2n2gz9
Swq4BBxZr6f/DkE4CXv4gaABRY1TB1qMxgTBh4+rbIcBqBDcXKcILGW8ylQcGZ2RuxN/xVqdcRNo
SROfiA65UyhacHFtRufCj4o9Z/CrYLsjGmzG82qrealVyV9FVzUYgMpy4M5O60jUvfc0S9njIFAP
QcZJyyURLwmNS5u1toVRVIeasGBM7mW5ry5w7dsMTU13U5sQCgD0e4es/C09fihIlqaqAZ8agOG0
dMw8EcuZf/Jcm0FtabdO1RVkWPYrAg6PlUveYpXba0KLxshVrGMenPE5EL+0bseP3lzotVXq8SDj
Ig0gD39QgMAq4e2yRWuZAphORaxOLiRHxMLQ43LtVKV0cF1eikGbwTZmQAcC+j7pzJRgfRZaj8OJ
v7ywKNatEktza4BHySlB6WTmVqNTtfnavoMUWrUvLhT4+ZP+qvGPHyRCHlVZDdQT0CbvipOuHG+V
cFMnq8exfFfH4necGY42DVvzjuXbL9/WfNggdVCRR0OC8EiUeXcpllk9dXheg0GK6JoglDGJNicI
6pqRrbv4BlNbMRJxlDIOhhKATNfxMiPN441ssi0xFNC1xiJ44JJBGZBeWPZiuDCSKm6FoRannwr8
viSFnlU9fpxYTvJpM9UR+uDi46doKE2hRsbYzVdbrCGjE+LjGkHoRBMPUMwbgJnVSo2sRzM4XJt9
AX1KmQHY19FRpAP+IDTACAyTvMlSdK+qURh3GHEbSqRPFA2paX8rgjxRcJzVAb1l70c/roiQms+x
kmaqd98mrhUArg287ucakpynzKyjUDiTYC/oeUIn1VOuB8bCLIq/JmetSy/s5M3MqILuU+Qa7qOW
7zK5Y8w+0rV9tqYd7WWID0AXrwbGmSOO0RziYH1nQ4obp/pyhnrhCAQeflmHxGUZu0Xa5KRfzdmx
FAIV6z+6tqw0ZKUZ1Z5zir8frzUvgiINCpZAoLbgMb4zIwCNLLueL4pYKX0x8ph2/JJE58hpobny
wFZRGFtQF8kKd6BJgMRhM6nznsmh7opTNbCzluf0GYkD7OaTF1CbxSggPzI3C71BS/8NDV00FxhA
4FmVC9Wt0PJP25ZaMYZ7dWGftqbbdeEaznAZCcO/jXUnEtGcrqwibXOD6BCpNjMARsuoVSa3mO1S
Tny4GwVJm1KrjJfGKjf1ojki2D4tTtthbhLhzECCky+rbU2cVYrWXMUElgXBYcTNgrrbSnhwJrA2
8rYCr9XwiRnh68oDq44b1DRi/Xbhisw0j+cOx01OTzumc4qP73p8lJC+87MZyz7XUnE8UiXzlsc6
bkWOj5EwtIIQzh3UxQ40nBT2ce2yKI6sPA/0WvZqFsNTtFAb9S+TQ8ZZ96InUJv2uwN5aViMDgtW
2ZkrNVMiEtQVp0uukdkWH+M3CwmD1v7Bei0afHbqvRn/SxkDibVYWNspPRuCeCQo4mjZRG9Du2qQ
kqzT6Ea6x8tSjsTwyY+jTjFe5O87lAy96neAyI3Iarje6yQ+QHI0QzLRlWeTVQY9s7LqLa7+zwTk
8kx3gWNUshqMxcM0WIGykvl6L9LpAgTwCNlhZvQWYeCDVUATtXyk/flTSDlNmB+/Ax78buifN97j
wYxva2Yu5QejowpNnqpkjpoLLGziZkf88+w9R/Xhm5ys+VfKhKEgD+gmxEOLCkRpFc0CkmI1T271
l3UYidyjWOXoAZw5ANOL0iiurFkLuIqzBAQAQYXPQdmUP5YZLOvm4B8B05kqLcI4dbjKAOJ34VUX
JDOn838agjO2dAsX57loZxNbaVKmHxQdHeRYJd7VcxRIxZGF5fqxX1PUu+8urScdXv6nDU0QJ6Fu
i1txYwblmlmkGnHLG6BgtxAjKbXO/EY5+TfaNgBPXSdXaYlYLlXv6SURzVe1GzOH8O9ZdXdVStxf
mmls1WVimgYhEJFTP8yyI+ChJSwhymnMXDJH3wx0stCZb4LT8Jl/g3p9KSo+Wepy9SC6Kn9n9cAa
A/FEoydIOmK1B/QY1BiRhbcqLsPjUSlvMmHVekBHVO4GT4RUEPIQRslPicrS+RuOUGMSk4+VKYWE
E5nk0EjVdDQnpLpyApmRuOaYR+Y4Fcu2qBFJvSnGlpUS/6z44LwGYmZe+qiY4RMiMtnlUHg41RJ/
thW9ckpoI33fFo8sD8mAquBhdkWlSYbcP3TsnO5N1wLNvM9OgMWmOxdK2BhRoKk0fEjQGoFeWJM+
YWjT2fdqoZz7iFFQT4WiQvHz0Svoxh1PYcBEWGGHfvqUN5A2rRdOQ8ur1U1qzICU08M6vZb9LeD2
/8XWWZm7BXSfAZbdVL2DP9EYIShwg9ZW1XedrT3+E3eJeJ8Cm+xaZv5rA4QNQJheKz9ePo91Qihn
qyuaabm3+52Zp2mJCYf8YHhbSvetMdeeF4UBTfhA/khcSGcqlDEsFXM+hx30WV0am4wwZFbxb3oZ
HuKzxmWemm8S/uwNAGRboQF45i0LPBBa+VPnYEeFzs7yWEq2caOJZKGgEF+gmQcuvF73Fc8BGv72
XMvGlWG3/O2Lup4qd7Mxgs3XBunMsWSYYmjxZqMEEzsYsgDIQ/cZ5Tv0nibkeJhlSXV+iFOUZbP5
muDj8Dqv64iuIFmT2wOPg2DUSty5YtNMB7OJ+eXn3/Dj2DXXT8XTdSty+H6bX6kdgXGhqAv6jsJr
76vNNb5jcBWIvG7to7iOHLe/YuQSPOEjEp38rQAaY1BlChoUsXgM2tbq4HOsE0LOVN6Lu4/bg6HQ
Wj9VoqLgljCsH33ZrgSoPBm3G5CB4fcqOX9wKapT5BiM5mu2Yjw5Wtq75A877eNtaWO7xiCIROL9
knmgDgGnDJgFytINbmR71mf+p+mf7S4P7w7gmSKBhjTOAFGr5hxIwJh0SEarGBlgMUlSVu8OiqFQ
qrO7PsGn1+/gAhCm9KmUyJcltnw4vr3ivtAIEQFGmFKNzGDDCIgDrGKFlgGvY94kereky05oOIfq
xIbipqOBZXDO40OipW03JRu1hblexqPNFPuv4bgnGW7Kb3Gbxut0MycPuH8DALFkKtiRXf7ch+hl
wQb6W/1NC1KTobdCQSWt4kGsbWdAXNbMJxzZqUjP/tMAiSPSZY8GRhRJbrDgjXsEAELaSLOpradd
mohjh5wfdmMlBtjlsNQb9BGS3DwqoXAUj+QeC3GzxSTqLcyfeM3DMDe8EFn85j05KcMlU+QsVzDc
xn+yfcKXTKF/Rdmh/PSbscta4RgPzNQuzAYbssSBskhaMWkhAAbXTT9hgUfIoQMRJuuvQ2SJBuox
dRhKpsKqBIjz2fdI1XX2zjvo5GpWo0JVwAEcOeKMwQkjtKavMdJwTkn9ZByoblvCUnPvNxRFOBio
UUjA4snmhAnEba8WPJuT2yQOWPqZ+B9edUxAnGMhqhGyHRyFGhSl4h73Nh3VhmvSfGX9iFnjEwdy
2qYEyOw9ER3ytrLxuXsoSgqH5ELKp5sZTB4FgXKko/fpp7mai2vLl42Nrvd6Y/NsFFQS2yWd/Bzk
NLxNe+h726kHr+sUweeJ6WB/RTG+gGqaD9y6dqlxXd6UnvZzHMBnVtAF0gRD4v3hwILWPdbm42FJ
/D7DcatPD6rpXuOBntJgGq7S38jlxfQvtFBpno7l9vInFUU/T9fQbqA2+cr6eyIbSkl6MVdp/a7y
jCF6/iUQNB27ZUrf/vtJuGY8UuVaMNgc9OqZFpFsEmxaUe0vjbiUzfxcGqi7/6cNFArmS+mWnCZW
9rYMNlsIUt43aokNu1dM1rvjSLYLb6S70c0rc7038MG/YonN2F1kFr7+eP9vytKqfUktMeWD4Oeb
kP5RVsSqzBenP3MqW8qoumjr3qLltpprfaYo+J/jNb5Twiy2XjVP5g1tQuF/EpD28PrNmeJFzOTF
mv6WFtbLnImpAMVnUIlzeGvNCJlrn8ziSH6qiTS8dSlkz+zXlg9U8oUPYrXJkMZmu3Sbayx2obKx
R4Wy9rMWGXMrMqzxmLPD59TZCukXaEooLILRyxnxXxMtFXB5r8Q3sS/wyUY5lMdcV3S8mlS76gNf
ddgndtv51SEtKqAraXiwMMBk2Hj91aGMTKvQja+qv9mvCk2uQWb29g1/Ypj93G/ofJ7igO5kbm2d
EeRtv7pKvBdh9pHz/b+vvP8lsQIFULnd6FsubtXDUW+EW2tTw5ZYKZLguBNrg+BMCoPfEMM629uh
7d2WGxfeBohPlOtiIEC5bolrCmIjud+W/IuLHgE8Jl3WbILn/4gBwtwXUc7e/2BLPEPlJImSigUu
BLoNCvBBcE3T4ZLUL2X3NDl5Qc9A93avVv8XWL4AcsegUfMn3b/zFaRDjVzfGJDiUyiJvnGfWz6T
a2lqagiKf313ChbKEF8wDZde8bi2jGhU5qDe43dJAHKgQOZ6RuGlQ1CxOU4kvf52HkM8TyUsBNDE
bVGQRW2Qh5TRcK8RvUaKgE+4ZzvFdOv4FZslQZ4ZfZyfy+CFwJXBWYMYdWDIzoKVagjMtKRB8k3I
kNtd+NwpB/XPo9RPU+cWp8NwbOdf370Z2JSfnHdwGnAzImpWPKlfEeffDgOpNmpad7Dd//qyXhsl
dV/jaYT2s1jcTh//RAPCIcdkTi3HSArq0pXOL2K6vpxI5eufhsFZ62wJeXYh27s5oAF18Hgd2URO
LfWzbWVqWuvNta3RxOoo5jipfDw+pIzeZFokLDcAVkNzpBlw7aNZK/9UFF1qRumW2SOo4lR3scel
Otugu9bUOHHd1HUdnHbpDkHqV6XETehehvZTXZtKQ9AoW7UrWL0KgM4l1BH3akTUtATzgW7toHVV
umYd2YQACEuuHqkWZ5HiDpNgtS/NlIRuZGfby+oer7IgpqbY/pdnFmhIlOib+QzntMOeMT0M21UQ
3QhNATZXNru8RhvGa5oUFYiSv610+6g0N2oA8hkAEs0LlOScH80kIP+LURPwfw8wqL78vMUD5g4s
o8v+IU/F7ZCiTxJPQKuSGOHDrLe/ROhHvEFwcGro82XTdpo8vS4447D5mfxt2RJjRzCgGx+1aZuI
tTGgUY1uFFKk8ESHyVRugOc9KnXK3oGZ9mZfuLbI0WI2ySZxcj3tbIb0y2XUj6Gt6KChEatiUTrW
KuQyXwVYjNDcPu96/eUrRiX8GHUDe+jezOtvDGjLIKY1m0KyaTe5F+7659cCj7DfBi+w6jhslW4g
Q/Cbzmh5FoddLRJkU8nOeMH3L+WecYaDlkGVGOfNZEh6J6bV5RHALeieMBlpoFQFD+At5dSrjSMb
DAlYyggoprLHrnLrUuC+T8NtveFbfVUaLZnQejbeSMX+0erYqcCYEup1R6NFxWf9LmW8OGWElkG0
plu5pshRRobSru+y12SCaaUF7PNSCfDfETAXe/efc7yLCfFQztTLhCUqscV8b32r4XOB6CITtQHE
s1I1pNZu7W6+tqpGGvgOJ/TXffjrU2IpdujHjzE9dquQ3HxbdZtwuZN6nWSZieoExOHe0aWuqym0
aTBs1v1tqQwfbDriDaAWZOLvOs7g8Y0+fDKSeOTWF78qg5Nj17yT2go6rOThcQlhCvUeaQUDDY6Z
ZZhEXv8nghbfDh4VtaTiHecz62PjXUi1E3FY6OPguOWlBs/UqHSYaZP2/sL+19e0I8o52GgXi0kW
vfEB7PWoCbRXBp+JFLRfzIDlx+eT2+lPo6MhX/tpCrhoPufTU5YetQYhNFN3NUToPW6M4kCpzpDo
PT4FZsaoCthDm0zXbJ2v2CKxkvoXDxNpIc66Zk9/Vj+C7Bqa1Wx4+JvVNuNFilr5Do1ijyOZeO1Y
/Ek8ITnwlDzzm7Vsq0yzFROYyDCqmZCiCygJS5LhCP6cHfzT1a0V/bISLQihSS8z3yOOwRZh3/rr
Kc0YuatPlaP9BIzdJ6l7Vndvlfr7eadcXT/xBezHgqxyPl02Ed/Wz34LBy3tcfhSCWctdstbFxkX
OWAAjFiAiCKpq8PC9C3+dE3RmuxRhOHsyLc8yrlpJ1es215X9qv+CiQWS2LY7/eHhzwb1ujRuuwC
LHlMiS4qEZpVOZuC/M5OO2rz3ZyTHOxLqrKQIIk0g5wMt+KlE4ZpvBr8oY9jsexpRFT3hpjGkJDi
okLmdWpVAVxI7HdhFdXb1lHeZEZBc8PbmUwIshh3gGIKI5A+OcxRD10ze7l4Pfkg8C8qpFsjJyiV
frIO8R6b/ZqNFG1G74ZWhyE4FNA8FPG/Bf2CzFgK+9RjjDSgrjBtyF+m2BvYzS2+Is2V2krkNp8z
DbOhpd4tQYWmg3kXS/mQNou/hU6UiuNk+DrWnBlFSBLaHJelX4+R/dk5dhcVHgiNGlCP1nUXPgMh
y6vM6DYm1mC1F6SyXHsldhmjXCAehnaknpvhg00qh9tWrPxc1Y7jIUCLDKGV/seh1DmvsdPfVhzs
cNSb5r3h6LV5tsHt27lfTXLSestaVStlTwjjBybgUxP2blqpDhlRRSeO0C26V2xFisDhATZEV2Fu
y1McuiEVvTRbjb3Z9K8fo+cKxbNBUY9AE9okKhdIaJby2uqYZtzOtoY6B8x3ea5I02XZYsjAkdK3
6XOcNzeeiirP7nGhbuYmqalpnz1qsm3lPO7I+BoOx4lQYo+M/c6U7cB+j6Ms+ei8FA4ziYJef6k6
sZAz49GNfcyHcccb0SEzUxx/DtVg1m8qSyUUmCFkWB6jnt6+IInFNIqh2a2pVD/edfkPSz4AefOw
jQUBSAOYBx7Qa4BQf024z/pwM+8eQpeqskZoFXqKo+fgLRBf+Ve9RT10lwRbnT5VTcwXPl1vGCzJ
IewcpIulYGV8ndc9eODC2VOzjqTtVE8iRuD6L76rToZlAfTNCqAB4LEus/MJWrq2bRyLDZbGGeVA
MPCpgOEqABHzLP9wtNeTBBPcDMSDHy3XJ8wCA4xOCTkOxhs/liUCkBbk8sRvuZLQVxX6CszwAG9c
3220Odav9qWKtGErNiyNabW+vZTJwyXhA0psf0WvFoslFWmmvsNQSCgh350YsKgI7MRfC1w4phAo
9k8GOk3NehK9wx2RK/wO1tJ7+fAKYvZSQzlUSW4CN2uW9AJ+yR7+oLsh0kElgccDBlybMRQxlU5g
YpOXb1v9tU0tp+Kcc8mFsLFYMOVVtIQnz13GN72CtID+bzEtKznN5xMbP9sBYl5+xene2uUbytwZ
OnpTm5PvhzvhHz5UTJEQjs1pQeWJuJSZQ2XyQ479YyXInnN52/MXrZZiFUoOdX8WM3oSgH4wY2JK
lOx3YYcnu8OhsLrm0XseUcApx4KZxHW/2xQscXzC7mh+UgdPoChrGdns0G4DrSCqFlhirrhCp4iM
nvFMVksC0SqB8uxFl9Bryy70beBl1w/AKbDTyQr3vM6ItK+c+JykFT9Pd2iZ76O6HflMbp3nJJ+P
ZosYHNlDcxWCXUlEMJT0mt4jWPKT0Uqu/LMBAUyGJ6wefiY9KuI1x5ks+IY1Xl/zAxMuSw6WhKNQ
hvLahN6AuBvG+oYQKRoD0ZEC2EqSxqdYxjmZBXlk8BA0BWkm3sdLSqMnamEYWRw892tsOzgFOmgl
FKE4/5C9irmiRP+173i23Hj4hG5/1Ya6Ro/f2SkcFLtyKzu5+Mm0XatIto3KltfgAF1mQLQwOPU9
eSVuIoU+ifHapJSfg9hg5C9D/5W6nebnQ6VycqMzB4cgJmW1L1l/9bMYSVEMCMFGTGv7dgV/4MVO
e0Oq7l4uW44VCVJ6ZFNBsa1KIfO03y2sHZ8aLdyRGePQMmXk/itCPMrZvUEIelELPmMzyXM67c7X
sWzPEopeZ6V3t9JVDdk7c4ol0U4iF3E5LMTjY1ZD3z0jBXX9SvSwzsazFMKlkjJJlSQYOY3Mj0sK
C4KojyD6INwd486Cy33YxKz5Lg2avNLuhmvd6LeDGZ8XdedDmP5HE8bw2sDCXkbXJGD67ZruhYXj
wBrMuBfNGpWXmlknW2CNbhG0nXi/StOI7B4a3wr38D6cY2Y0GOYYmIXu+UtrBJO+1PMZO6Ni2dOl
JBG9yk7QHY+XY1FYZjMVTY+33GvTDTjOtWTTskv+Yvk4BZT+U3V/IsSsX7A4XYLpq5dj3wJyY2G5
VCP/zcOQe7sVDeqP7eSPA7RF082ETbZs4sc3meQ5FzmDkIocKq+NkQuBM0ZPDezQTiNisi8NdT/5
omwHV3fiTARJz1VcWIpQug1T3c0xCr15c7Kns1QdBKONz7duYSkdvHFX+PA/mU9Ju9vexLMhjtFY
HhcQALrkgR5R1zJJ4XB/I+6npwmreB7cH5SoykwOltzia6tWkYEV0adeO9I/Mjh5VntOOdq4bocZ
AAC5GpgFSJdsQtfG1pIZDAMyu44gpxFgYkavX9Yk3UF78jLTaWV75rd9riWmxx1I5fAJaqsbdYuh
q0MaDEFL7nceiX7iFedbZQ37pR2aAEnuQv1OqoDsu5VmIKLqBL7KOqA6vPrIEVv4pNU2nNindTUo
i4Qy8/OmUNAh+sdvoeXYKvmAz0+fqH2IejN74MnuodFCwRBNeAP8rBFzxQkPHYlE9vfKDgyW6cvU
qZKG6AohMq4dCYBm5S2NssrXDk0TdVB3tzkEyh9DvnhlnRySMHl5tKe2noj2DeMKBbG6K9GWzqUa
cAyADXkgLQgXmuOsan2pt0W1Yw13AGUgXyJN/+pbRyDmZPhg0sTR/uUuQBGigSd01GxlNjZOSnhC
QD1gH/Pd1WpUHoSbel37qkm/mpNAOCc7Pa1u03QPeZEWhz964NFwI0JaGhg1Smlsc2efTOBq3L73
laVG3Vd9fo2NFwcyG1+zXN4jBmGaO3Ybm6N/g3GcTy1h3W5vvm7oXIJFGhSzyHQXUO6TfihTBfma
bfiDuGBs/pwK/bJ9KfouweerszaiZDtWlfXQTf0mF0DBm6l45tGVVpEiwWHu173dhdq89fr/mbhT
hgE3r+LlHat+hOuPDb8wPJdTHemFe1Lg0HI0s/JFZLw7eZD6ena0pu5/7uxPOFxU5/e6NxN00R9A
kmsmt/pxu4Tt4K8d4+vld6CXUmSYNgoo4u6Cd2Q1u66np+5TFSYTkzieLbaUC9gpB2qTxRGlznry
3p3SHdWYJVbA3Qx+r4qCVTqcOnbozBouAEQKKpWc+rRwC8aP0W2Uf8NVFGrr/9fGNK7UFBbS32Hw
ren3XiDxGtKrHFlKbd06O3CBDwGI69dGXAAYpIYnORaLSvPcwcaLYXWop4qnlPoZoCwROUb8IQTG
emisoAMPrvaRqta7UeG9BocR/YomStDei/XUrf2lFdQwCK61nXT5hbSCnwKNECS9K1ZQJdj2KGh/
DDVxdeG90PZ2MyvDWrFR8a5Q5MLwjI7Z7fNc944lmb0Mfi6dG+8eMBl4s2ILGTNfGEqYqHh3OpA+
amodclo8m30OpjoIqmZL6CXYcJ4s730avgZRaQIADH37MfNToSkTAPlyEnZMa4q5cwettAv9klhG
Q8DB0t2y8TqPxq3zpeq7/YruZaZVCezKOqCQC+aHgyh/ajtX5JlXQJwuWGVTPnW+gXlyeG/YjSts
gjKsH1k96l/amhzjbVRKvmzoBVGE1QnHHffdyReBhNbaZuc2Q4MqTKbf5+DobYN47gbjQvyHw86z
1FHZqepTBANncriroZQkqrcINtbP7Hoh5rR5sE/aWQRWtQz1rQ3HWBIFX63/M+mWbk699a9BJtRF
bFTlEfAKhmJjjMFSmnyAIOvxbQCKtQ2EQgIrvYeKySUlO+GjhBrZeL0yWoPSM8Nops+4c3D8H2Fn
wWvIE/uaIXIqHkgeFFJYigeOuh8Z6HTSjErvv0n2qHVd2hxKSwMFaGEW/PiI/kpNydUs79TjZMJK
9VPfT+eFnyZDWfuXrVBL2ysOQtFH1v5nMPcTUimsSYrAXdnE329k4OKZukRJKQp5ND+iwPRM0sEL
u51Ii4S+bvnZMIEiPq4fb1cnkBeR/LSC588xTtJRPOnVJSYpOhgQ/d0nb53fSlT/xe6ZQcRhERPK
q0ngU55nOgbRdJUtUaiW/SfI7GCqiXjfDGF24jgMhJBgjoqFc+VuaKo+gR3M/3r3XU2BKDuabZAi
W6wF22EcWhPHaewVakd9b0tqYS/Dy+F1UZTagzfkepSkBuTP5cKL4F1MIddcNiuTMWiCyRqI5BJO
5zai3RDz4UdSsg78GB09M31Im1AhT16KpCLiCjnk6hFaPzAClD8LX8f7cP+55gRkh3cBRiMONnxH
NVju6KUekFiVP3jKU7wf0J2gUHlR9SbvzvzNEiTnNdETZQg+K/a5hcSjxMLp6HAQzAMbZprAEFYG
2fmqBDOlc7kfc2A2MhBW39ZQDja8HTUiEuo40kUGlNL9MsP55NfeTDukSQERrdUpypkEFaS7Do2s
B9gNuOyguK/Jg2UPqlPeegydnKT1QpesZBSvhQME2iolC4GK8SAR4dtkegFuxziFFyseykYLOBdQ
hRQflx2epEa5LP9SjPj1oydcRzXKKBrW9N6b6jEGV4z2Krz6FV9AV3F5B/hyYxCEDJygclfsxG1q
nDpCEhazldgF7UfH1rxjcb5YLA0rFRWPddHUru1Vsga8IxaIVT+JaMaOGR+ti/inBNnr8OKlNr6Q
ayi24tp8xR2cS5xAMO2LCTZu8go4K97T6lPfZLZOTEqcTufregxIr4QSI7muHhiZ9jBtLf0ZcSZb
EdHrIIqO+xhLORd9viQMbgHDuuXS8T6byNLArvy60emK+g8Gn9bT8w6xBfFh21kMj5EU2qoLxnx2
ymI4l3l6bAb+fd8nybwPQnucgojrKP/Bod04VXPvYR0WgZF2Xtu+c+74aowp+haCOoX6T4eyjN1H
cUtNdMUiR8y6zIOi6fNlM5gTF8m6mpzGEY723PEVmxAS8et6gJn81IUxQDBzXjnXvDn2bJzjduAG
V3vj1O/JrVcIVlvJzUIPtuINJhsdgKMef7/3aVvtLmhHgC735UKOgu5IwzeNLuEmSGkULL03rm2h
INdFbmvPmNCK6WUanHzvXba5LIzXuLl3jf2li7EK/4vdC26HMrKOJXRLzVHuD2dtdV69lyl85k2/
JngSAFlzUKrgL9i+ZCm+HnqatU+uIMNRR4Hscd+P5+EVWA8DuTddXmfdwMjUO3MVJMV4VBWpWIpF
5XJYSx67wurBYg0wlZs+ubOtSET7et+2aZgj7v7QgnqnHeHysBDwinukI882HPfRNgmZxQTTLIbD
iYOWRo8crmxvTRADvsNvnLs8fQCLi82Y04c3LtpmYf0o7Ly9ISS9sckqLK9IJg+1lF+q93MjcgU6
6PD1lLLJkmTLiJNyiHjT1rfHt1D/PUm+Db7W6pH5lJ79mrqvXkVn1gcrgGBXowyZ2R1lnEy6wUt3
SShxwx1swnT4deyx/vFM8AVjcziuT8sR1d58WuFkIlMtT4GGlCae1qN5N3LwHkl0fvJEH1MXqK9C
YjS1BzGLP3JYpC5IrpEDw7E312VSoHobuPS3rMoTxHmucT+EuVKrthBPVX6H1sEO297xeXr7hn98
EezZIy2i5NDhoqozJ3RI6aztOAMxe4LCrIHXYKJfiE/5+oqUrUtQLgLImudIa2VgOk16tm86JqEf
O7eDAzCgDc6ocMdR+C2KA+WsKuc44gPuM2HXVAr2ZkrLxgUHnYVgr+oTY0AXiwNWK8UAjkR3Ih7p
en9FzR6SqaOc6ScHzcEn1zS1q+Y7S8xfFRnH0oMXv8aaWy97N3YrJa3iP0xRk4GH0y7K81JWeAPB
CVhQN9iay1TAkK5RVw6s77ZGjKBppORnHkCAbjv+hK6b9XmiGKv15aAGhUZDtBPxsL02M5JklFxi
RzNuYYjV9hJhBIWUcFKvCDrXWBDH/VE6psQ7vmszcWIAJXJlfI1bmRXsfDmV92F+DwPee3KVvQ3I
J0SouapwqoYaoB4ar/SQJ6+TsIPYMqae6eOOT1FyFjv/CJeorw30H+s6z2b2pp0Mft7Mp1zvkn3U
o97Fc5WXucnUWdL6URkAmnp2sm77QxX6SPPwXnVeciLk7QHyVUXs30T5hx1DGPXAf1T7ouHkuMyf
EPec1dpxik3QjGX/REoJZZRE0LeA5PmYIIZWUN0CAEdSUZApXB6o3U9pXERUx1YqP1zQFNaLIWZs
8bn7aJc2+p4rm0dF4KtM8vtYzxYZMEfgnVDuhuphZTFvuLTZkrYNHlynKCg9KDchvDa+gvSgk7ka
bhpcq/7irz838esn+kEHAE49zvr6kc6Qy/t2evld7VxgPg79WTj3jRvewOlDFLotxcRMsOgxaahW
6pOhp71vyxx1dOYB6EcKIFSMOrMoOyPQ2zJvLsQucVWUnfu/QICXB0e7rgQImh9Vsnj1iROZulwh
g1YHcOmgjiwLkP0Bb5JOoWWU6fkL4pnwRaOMOhtVZ+dIbR+tZF3M0ErGYylUeGQjKqHVuXeKhOck
Q1UGGEU5VhbGcBRg5OoRJKfxTb4G/u5CtQStnKQHPn5tY6Bx+dPRe+OZo5YrYUsAg3rGfpzVFmv9
Ulv2hNSl0nSwMEtgQYp2HzviU1uVdGOsEyrpLI1brMaQHjHFwvS+C2riWqlTzzVPZX1F3jT0Xlkr
spvItRleIACpbGe1QJoK8MaqgcPFDq+8/uSBf/HkhQ30ZQ5RY+XPocQ8lYKkabp6Gr+Dq1C9QAeC
ST+/w02fyIR+mIjFAXgO60CdWjlYJnmiHGQt+8FY7UxgBx2DZs5j/DHs+3DjHMJ7xKsnIO/N08Mq
El2Yl7wZTBsZKNk8h0/Hvif94p/7wSIHegG+WrKMQKREXfpvW7njYBqX1K80/Xrx3VJLQ2FpsD+b
Xc5qRrs8tnszkqhuhJZXvxJw8UPucDyFM97sEe6zbSJ7pkDRwcwv1c2kl2yoyWa8EMOkerBOI3S/
vCDmxid7QKW5UeQikMpulq5X8UW3+WD5YapoPVdPLxwop374jtVQYxPA4Sl0JyaonrPcpdroigYe
6zMMPLi+swNhTZ7G0Z2P9n5m/l4DYcnUUmqQqLrGe20bMxQ4NIp1eijzaSFf8ocYefA4osaWCVBW
rTKFlzaBes55jDjFgw9HuteKBzIhH7H0AL/0cMQ7EvMDNCU1RQaezqHFKVXxXk7l0Ay1LDm3ViAY
qLj04VsNLZjqUQ2vnU5txg65nNMKe812LDqt1YvEOMp9rRoeWZS2J/0SjzPjlxThtpCyWYWudMb8
YwHEw+U6uND3hg/RrHL1Zc1+GhRBIWZVJj++b6SUJRusowt5MpQSHG0Rio+Y/ZioJdm+1QqNuhHD
1igHYeJBgW1+tNI56YqkP6Cr4us7gf4lfirWtg4hBubLYG5DY7Cc+sSjt5tXmPbmsE1jvWOiF6O0
fAxPkyKhXoA4ga8l6neuJjSS+++gfmUgncI91wFhR7RrRAKGyH3+QRCXRlzzOtOUcY178nbB/Qhg
RTyca4pd2NwBmOpy31/mlgfph/+WU3oyBn/4aZY/EWEflRGQxRej626Tc1NuHRN6YESNRQMZuZs7
QtWAWZSVvEwfdGcLsyzi2ghvBlw+KtjtC537KA4ppSMks64lt8AFNz2o2ziWvjSMO1jSYKeoukF5
D8OsQh6CPF4ZXhlElWTrnYN/SxBljRPZnWglUAsjN52FduAxUq7Y6NrVBnbHQ/dm6vz8VMRrF3wN
ZERQxI1icHWkMbC+IYxcIpSRFovkeGkAGRpDuwNsgCvPp4NRE/iM04r4kfAldCEeyIOCpQLhyjJv
yFjATZeSNcVqplWb3SVmubG5vSY23s/QP20x3IEMuF3/ZKFL4qiBxH78odLH5A/qLgmW5s02UmZQ
o8msQPj2o3P/sG64qJnOsL4L+q7G7pYuyXv3x3IpG3mVtXwV/QmLVjctl/Fao2q8cBNb4DxrFNBm
yAJGuZfpJeLJM/5/hqm6Wmcxxuf6KHONQm1NEXuS2qqAQvEzg4/9y3uaKUeVxr15TjP71hgMS0Su
xYesn+OsvduEK0eVDW6L1mQ4X+NoItVJ5ncQuBFPxDXG5HVq2DiiZ1biadHIwL6LYqNesJenw61e
stL5qUBsSSFyiQut/DuVbt0+NLgKCm6ounGi1z3OZKnuFg15AbSXHSlxcNgNn0Dfb74a0+0sqZDX
2vu4HqJ2B7mFZGBsrKQ4CeUgcFgIbOz2GGuVm3Orw4zreT2+sSerXjSUepJ1ekAV04JVU1WwTfiA
mpTEwHNglhp6kIV+egBVcg59lER95544Huyl8iVcAtj6KOqB0SBbDg4BKP0829NGtrn3n9ayysEK
/nrqgaKhPFXWgegAaykGpDqTn7XgZPHzUvOIK+Wd2ioUBj663Xf5r4t2paYKF1sYuQLlbgCbc6Kz
Jd/epmyCbPX1oF25Cwl2aHSHuG+5bqlpp7Cw4zJRow3Ql/63wdvsWr2UE3e+xWXAmtqtxt6A0iS9
Ot8zZY1N8rFNXNAgAmJZkKzTDVZ9bOH3x0pf+nXh4909n4hh0pNhpSo/lBWU2Qkcht5uldXor4Xv
vWGSd5ah2OSKCi8pf5spTp+/DpufRO8BvrIPX7eD+lzvQpByPdW0Ex7XoY1h+72TjXyZafmUHuNR
Yxa1KdwTKFC+3tB8rS0fMNOiDC1/gZQSq9NuxwWljxrV9SR8IxKXmZ7cbBESCpPjYSV+gHcvrJGG
DN0N19YOHbKHp4/D6w2wY5oFfMQuRDCRrlxz2caHRj/RPI9riGgIMXjWkJl9X9Ot7702UIOZ82ZJ
EQ7HK7duU53jrzkk0Af6eM1YTCHD+8vXN1NyJoskxJ/vlCOcvyAxIkFdf8wzcueetCGKnUwjWPpf
/Dj06sQ5tnw53EhbndM7K6PCiii1EpEb8S71LSZlvm9SUWBeCkj1yaPgyl9eyD3vyDKT4K9DWI4O
t5ZHsXCkOGeWtd6YJb7IPm2jD38yfZr5xkgals4MQOvMTRV30DFAvho99lyM43ahDngwM4gTYohO
dJ4XegWOwx3SSf7ED+FfJMu5auA16+dOqgSwJZlBrxH8EPFHaGBRZi3ay1BhI7vUE8YzpQmqbhck
6KCLiai7+vEguoTQGP5MbJRCT/33F1c+ZZovOKk+k8uyvMkN9KDWhPE4T9qHdIRTsXVwfNxAsV3k
b2J//bS3rX2fo/tbAwWe39jrrpaQ0fu6B5VcJsKfGR26dyG2jROwSsOKYzR5knK0DoVoE5qvT/iB
SXr0w8W/lsemNk2HDaYixNO+ty6FiPlUDTS+Eof2LhAQo4iBmZmsFEiva4cY4J1StTFsouaYNB3R
wetFbgYExwlcQSSkpG7i5t2Fz3DRlX1844f9mXIiG9Y58CntrdOWbZoN27MCU43lpFZJaneABy2N
yor8lE4rLvQS4wpOAT25kRgZs9Xe95d/kFadtwMYpGjrHESrjQEK7yN++cwJ4ep9v4yksk7/HJi7
g9aXN31jDQQrcV+qDNLpVpl4ue1nkjHAhAJwD9ZLI9NwdRsU90t5AWspiRpc3nC19vQ36NNPKa83
2askC613AicMhG36tKSE+X3aaQI7UqQoLAnFC/GU0Dv7wXBck1zuJMbqVkP/V6GaRGB2ogfgDb2D
LOs3vExvw14Ca4JDNORKKS7ik0znFGm86bCPQS/TidOK2rlrGcKGnjaxiuIM2esttA3s5RV73h9Q
WehJkxcxsy1M0BoiLBWpFikItV6sGNn4PGvzihZwLvdENxSUfinNuoltBwF6CE/MbRKhJVWtVuZu
b5zafQH74Mq7oq8dwi2A7ekKBoBs5H6yXHrNOjVew4RCG4Dg46KDK0cIK5G+KNJq8p5maGvkLUJc
MRF+8K3Zhen02U5QPrRv+WQ4iLn2M0pg0wvZd+uMcxSbkYrZ9igvdCNrP1K+f+NclhLcLbQm4xRC
qK1jWRi0F/eDwDpBBWvmmNE/4mge9vvuBK+8GJL5pexomPpPdeUD0os+vlKxeOLY0TSpn56MziCJ
bVxUsK/KlmCcTvrikyXlUwWZZk7gTsRRYCtTR0lomCGOuTN/8DccwKa+3pUR/V7W21p6/BWmt1l/
OXx7DUKRiIZX/b8gdmtH4OaSp5NlM4JfD8tNc+3VA0RXmL6W1fLyn+UShMqRwj3saMbt6VoTVF0i
TAzbO606+xltiB1F9/6IntHivlJ8aAXFTN0SgbkxQipyKaWGV0G6rR35YIwfuhhsIl6lSJJPypfp
7k9y7+DsOY9I6f91jyPW40qEv7Y/V718D5I961pkHRmeBV4KuxnDgW4zduDcr1FvsItWbD+7cb3M
iKCMEdIrT+cRH5FYkFw61BLnAvFpSh5NEQIvyu44eqi95X+nlwL4eOncxSS31XpRg8MaI/mf9Ijm
SVehEKpoTJFAVoA+Q/7MlJZmt97zqnhfbozoZ4lftYzp3yjnKnocUJRoeHnUICsl0Av3UwJ4qbLO
JOM7p+wCSNXtfFnfoUoq2mn/f0f0BnRZ4ZSUOm4UKCToksEgsuNYHxOmFsyUsqjeUguP+ujn4ifT
J7WyNtntjZnT8vcPgtZd6p8c+C30CDn+Gs94A/5Qo+7QWPzbNioXndFzoghruHYsywU7jysScxvB
7XvYZJM86dt+Mh0VjhUAptlyAVXr7piNalbd/k57V2JCGp+hvO3enBi0AJ5OZNIRqBWVyT7sDtDq
FUcvtZWK1w2NPbO6by3R8zYgz3pD7cGyg2avbiOrI/x7DzTxCDwECm1sPfrfFzceT08mRqyvjGaC
+vvJ5u9Z3i/EvedJBQ2H/LmFNCfwcLdBVIgsHn3N2qXJAtjkh8lT7TAfrtLir27g7oEONSnQFj+P
E4ilCErfUOelMUevNDdI99hC+oAMZEmVLV22mkZdjKJUl93BRwSg6eH9RD/tAoKSJqDbbNtSrjZV
QZqBZr4wKMwO/sG0A0nBBrHOVaz+64zpJF3f47hwuai2yGTwTy7vGnbfeSzl/MV7Gz1qsL8lBE1M
OIpIF4OPJtssr7QDHkJM7PtRW0ZQgLWMVNlBTjqDV39fGTsFhrMv3Py9rAB1TYCHx2uiJmPEbqxB
wAacylunnA/9ZXOMNIW5Iz2UyNxfn303vF842wbSBJImZ5O6+XTbS+ZgXXJEp+CS+kCZ71hQ1i7R
a0lKGXcUF8U8Nd86RwntAIguAZ0oPK58ZoKtkmIExgpqxlPfVlMNMqnWn88UyiCizJmnUIKzeNJr
XLH4rw3SH9CL9U91e+kAsRVEcwWw/DJpRuSc0WugDH8CcHcVhp7DuiLvr1OJEWO4tSBBeju3VE0O
U44IYqGIfPbvdh8+tJjjnuFbvo6P1yIe99PjanrArtmKyMXlj+l1tL9MPTpXlfFaBlWj8BR/XfRP
9lVfdVZDDqDczP5Rk8to8EOdcbyV4pUN1sZlweWkVOwSIHyMMCGmyC/Uw48KPF/C9jz5CF9x0RrX
h6PB/Pomk0yvnxNZMqrZ5NFqA7xNv7n8fRxCRcuh/zNDzYxTKpBNTuTGa1DvFM00BsYwKClQIqHK
Euf+oJ3jvJct/A9tee8I9cDJRwrF+LLqTvu+rjZr72ukhP3bRxoeeMJQCIglu+SulOny0vMLywIo
rQFx8jisGSTPEgKzJNYD16sl8UQxA2S6VOVF/Svmz/LZDk34/V6jQneE8tCXRv9AgMfLneOEjTjc
u2X81d3kHE7LuAvNUP7LvMFdx1Jerz8zDDGhmwJKAF7dmVT8drXGt1JWAfl9Azx3W3/yjZc9pHGy
ir68EH7gbPBYRd7TheBqWlhR+GKkUoH0dDaqpktNPcgiLRhkjo1oyPPUTRQbVwWpAtj18fQCs6DO
j5HCsF866tsb2BDvB+bSqp7z+4T5YC52GDZHEuLca35cFirIrEHYn52lhfhM0acORhozNVSYpL9s
WLi5cPe16wR7lHdOvfJ6S9XPPfSGt8LTsfK9C26wbjqge+K6ZbWMzTewyzoZOYxTmy3IBEpcGRTo
54pwC8fD+FHSQDFvzYNDIXxpBKdaBC+bMG27P3+WyDCP6z61xlZRqK7KpRKl/Mx2PamM+YwA0J1y
p/jrBD7iDAdPEO75kFFDKGErQxtAFq+F10DDG7dKsM0cyH1KuR9sePEGA6rL4vjes0/CYhN5hxFL
t1fNmo74zpfDtqP31UYqjKA6EFU7aBLfQxVTtb55ygh9SGmHcFf4B8rL7IRoIs17IBF1Q1RtThHR
sy3z4i1uKtTk9f1gibAJthBYgXOWzK6aQYYfDC2w78CXFV/4qu0BdHJYQrsyRHkFe/6cTynOH0ny
bBsdH2W049QRpTwWQRzT1imOZCGTBuZb/ASrZbtgOLbJJ8Y11mrDEcej0PlI8LWA3DUAivmYWHdO
3CN4+d3PQVwg4DykphMoXsIoeYNnsMSS1gVw3f056gOzcnA0xWtMwlw9VmigP6Spmw0XDAmxHo5h
DnsBqzimR3vLO6Xk/JZ5riOVOjpBO9Tx3Rihcr3JB9EUW1kJUxtTBNx/c9L0mwCjOT7m/gTmdIyL
F1AadyfYu2VuPt5qzronkXSlnKcFLoVBaRmMxb3whjnJCsrvvVJI6oLwDWraYZBbF5TDAD3ooMah
kC2RyU8isuW9OiPCBzPNYgg6GVyvkPwhqCpj2VGGxkfrSD9hSFSr0Um8R92b8SEacKTdk99rfn/O
eDS8gCXZccQCBFJfrZzBRSAIPUaBHOBwY+zOy1leEMM/z/UZeEA+PZ90GB7aewv0rSFNBlOMzr2m
MRLQI5N0aq0PlKh1UlAJTmiLKgci0zTxAAXsjsAaCMclk9R24FA+y2UjAUoC2CztjldBShYC/xyX
VqVwTgNJXLXolvbqx8cF/yxmTEPJFDT59bdc0GJBSiY5FHQ8GgVOXQrcg5PePAnn8hTi+oJ2FFTm
8chwYng5DnmGx6I5tg0FNEiC8SP/3VswZ6W/nbYWcXUJntomNioo3tXFrnkj6Zoo1IGuhdcwQYAx
JZL7jR1144E7MOaxmTwGc3fTt1aC1qO7UyUkYxGDnydCwg1RGzEUn20DPn3sMXT6FineRRvXvihn
Ft1DK70YAyTG7jo54v6rN2GWkBPwZ+xWc2vr4H+aZEcyn+HgoY1a5wmBmjy/YZodwwGsaXGzcEli
IFUEIzI1ZPJRWsWv0bGOgUTk6E0vNjBR+1ZsOl4ykjJH2KRCP63NFzzQEUSLwB7V45OdWWmUsVuo
G7yyikfqL2Wh37lnMU3+TXa2DTGAvejvGWgCRiol3NuRAxnfzw+Pa+Wp2f7nVQZjyM3jvhRo17EH
y7mY2GLFh1aMY9mpBOUgHey+tlJx7cXudTCW0jLN1TNUZUa2z92JNd7YeuvsD2BIXQQk4kIr83y9
DXcamNbuvplbluaK1xfrpfFoLpmX67YGtHi4KVhIC+OcFpXcVpCuyN4oIZdhYvayz35x8h6Cs5zd
W8wUc5alROtM7noYqA+IJWsL7etgjs1Af5B8XwUbrLe5ck0UVRhuCJbQlHFuZv9QWZczTMXC474w
5DPdMPbJUAjDV3NDEM9s50swfJmPdmZ1cc2QMurblkFNrtZQ09QCzN5tl/2DJ4o0Ze1CtUI8a0UB
2wrVfHvkXU69qQJOlzsN7QzZJWSZnNSG4j4AkBCWX8IlAwcISFyQEb/oGm/QKL8zBa2XevpBUpuH
LGeq9F2zQ8oZn8uBWFb/gUjKdH4fYVQgHEH1OwR92a2RRmP4Gu+xJSAnuVXUoXEATPLzuEqjgnLp
poGApEQCJWOAgZU3zB7/EYVdGpPMw4lNkppeWhZHZcOPTA/YMWUt1rFbvcs0BdugQt3ZE+jl1ONx
mJn6m/mc06hiWk8NnxA2RAmxeySSMJ+gsYRPKdRkgqXqF40S8pveatiEWHxtfQv8V8P4INslekLo
C2DgMZ40edh+I5j6h+XHPKJ59aDCg+838SCGhzfaP92g3iNlSaXeUyd6AiebVdcHxx9bZH2aSFoH
U9fghw8FgyuFARWKzNwEsLRZAecZIMt/7HadHEqZGPXSJ6Ec+XYc1gTXjpeS3cD1hdOU1QnoK/tM
B/JltHVap/aLBpsfaCiYw+DskfgGUdpUJvkQfd//i5WwKC5BM4Ti+Ut6MqPcO/emJPpHUrYZcbD8
f82XEEi3dp18jCs32xcqTwPbX2i0JG7g0L0jJsplPCHiZL8HWpEPXmmPXSHECRLv7z7v/I3G6fiE
eNnPTIK+VbKIOVizYotfAncESBNXhMeUEFsUt+gs7asULt4hzYmUvekZEAXB6DqruJl1NI/K/C6R
jVfsV0DRWio1J25Fwbbf16O1p991JdBiv1QCHnzaaJly41AyrudLkwfoEa3nTwVk8Nh1IMywwRyY
/IpKiIQ5ZjUAqQz7AGlNWlswkmHnTFGW81i7b7dSpaqGypcP/mRp+ejcMwrWqxlJdookfaFj4hIk
UFU6c+9hacSi6DU8y+JJS1u0X4VLXFkCidGHQQLlpe1vi64ufe31vlGB3mXg5wRkgWJEOfIRgFwJ
JQS24QTyFCp5S3mU+TgoBWhQQrft9ZO5wgYb4l0aBKoslWGVIqj/piJfDtRNEKUZZwMKZf9CEskp
0/tOx7fS7iEZBEl1nDuxE8Z0vb8hJjqml/m5NuVUJKgL99WnwI+KJ1S0x/dfrMJEAgdn8DgPm4FE
6/P7bMa6XbCRBmxefWoJjx9SHqpyOpFZ9xDggKif/PXpPxLIz3mosW+ozeJmzQwwlo0P9Nqcmg2q
vMwdfzCeYAFcnL1uSd5NKfKcWFJatmlPiOebraRbcEr6KtkgD+Ug61s18lYGO777hea6MWP0WvzB
BgfjfOhl2/cuDS/R0AmT4VLYSCx+SXrzsWcltzFqx3PjOKrlZjWo0N0z7EenszQ0S0KiIX4ISzww
i+3RzioSYn2rBNERyYixLY8uos4yOigjJMoTpn4kW9RhJMfRcG3rkdkowsBY1Kdf1WHhtTYHUOrj
cjhIPKTU0Ex/62eRpY7P2R6l8ZVLn3S8J6c/tvZScNFvjeoW3KwWQ6mBkuu7pPAQ07xaNgYAVJoS
gMd5N2wDUJSOhD3rv9kKaRJM7NdJMuNFv4af5BFWzhM7HHaG7bOGoHEc5tBTbG7NdRk/dQ1bcngp
MrC23SiZ5Mbtq9ewd2eXla9IgzCYJssUWhinFpgijNB1IaQP9N0BEMADXRAwJVFtiO+y6tQUunu3
BUv+OTl4iEonMFA1DHpPzvfOyzHc0xHKS6fjB7wvPj4tGOm4jtuHb5P/kKNDfItR6WMs2ReEj7tp
wKiq4FFTYfqrYIRxbUVd1B2sjvUiqhYIrhU/BgOK1Fr9AcbDihdUU/oCiDv6AisGdGwtfC2gwi6X
40G/vT/7rbg+VvZ2cQwrm+lJ0LPIKrhzjRL+YqOf4klTeGZSKDLDdWl/VZ7wEfUy2c6rqXu3HLJ9
WjAG9TM6jODGjnm4sbUAM89Pv38MZ7INIK7Ib+UZvLy/DUz3tjUIvfsLJSJJeQwOP93UydB/NfjJ
WYm4GfI5IGkoyjVS2o6osgrvuCxiaolGD1HzQWMkqQtnCWDzxhlQ0iQp76x5Mp++fbWlp6ohe2Xn
R2/yjpX2cLHj7FUGuSI3h4vKOWlpRSIDuoMPCfkoT0kLLFbD8FHGZ1rE0JZJ91DrMpRF7oemO3we
jxjocl4/rwftM4C6gE2jPRkjeV/DckjLsM9vocnJs96pcqhez95ERo+KOoM1KoTfdBZ5d04gOkQQ
j2k4itlEAxQexApowcPScZBaybT7u0bjRNqVNT8YEHYoqTeoNxz7MKmg7+FaHMk89fTuLaXy2+cF
N4Nr0vGaq5btU4205OqA1XRdSw/ymHqvN/DL17jnbVR0eSWjLeqPp+87G9ZtL3YCKFFy6kIb2aIY
oAouJQtPld3h6UJh0XCqYSQ+BIM3U1067UhRPBNjBVVuH4a4KGmKcOVc8OJ2cIjY+1QYQ89SZ1Xh
JhZhhvUCBWjtvCJ3FrEKFAAnrC7DxpeWwyElyXKImMSVsmdSgwEuRySFgsD77pAgI/ZtTIr8+8Ak
I19i8SlayHgXyjeQXyTiOCKzdy68/u6iRHcsqAnyQLWZShbIjI/1GZSTST9q+QuWXhZAShdRGK6C
HCTJ2a2zLLxuEktqe3r1s7Au24JHKF18Gk+mapyGj2xablcXCi6/WjJsqCNyTvNfoE6gRFM/gASX
5g3yNJvz3y8FnHBkmPYObDL5t9VAzyam63nX0gJatnSbpAvfgsGSenr4KJyiVAUnq5zTFtVknlGp
hySJeOEHFTfw6wrtXHguGE0BaCAhWn1Yjk/2uQJK3ZtAULG1qz5w42CqJiC0GG7FN9m7j1nbHuck
RSdqMeykT/s2nzV9SzxzyYLMPEEk4xm5wOX5mcH19AWGYL+M3yTnwc8g3zkawRnP/vbfRUVCz7mE
Y+Q0bM4olCwSqTWlkaqw9I3H0P3RCbruI0BN0pJVrWySzJZksMRvnuycARx3bFh9fZ0/Zx03G5m6
tdu4GPmdaTQkD41gPbmPuz1TCDM+oU64DoNNtkZb9Xv7PIdK/9LOBiNyviRFBmJ4MCBkHBNudXAL
anLoJR7TaJSxPRW0Hgns1JlhSf5rIp3zXrFFTxT5UIYl9yj3SKSH9JGBjLy/hTwDlqqx3btp2MwO
p3esQPbZ7in4JZxoF7MwGMbZY68LmcrSRnVCp9/BuKy0ZK3jvaO5GMU++TsKZvuv3Bv/fkhRBsuq
+KQtiw8wMDMhLfGErCheRvp1ggF+5gzZHYcNiJGWlk5XcPu8hMVMuyg3ppmtuC0JcK8txtCcRjBQ
6ZW4kLEh6sghaC0tmEoP5zQzbW5QHL+z1Q6uZOsi3bcy5utkMrd89SU0NyiGpDbxa74AxKrE25SY
s3rWs31ATfGZ0TktDnCrWFeRpC2ItFcpQFcc4ubmnvQOOXhxmNi+qhXa4kEBqnmS+KdqQv0XKflA
tENSGLLivPoc4l0hk/Sc+9D+AFC6V6/6b5zVJ22CxS7aGX9dEcj/ymuCRZgsYzLThLn4R9ft/G7c
wP+wIYY+gAts7mM5cjWBGShdgqztoI8lVhwGkEvCI2hYKoU1HmAD77BdMCIpAeV0FGqonbkK9CNJ
eCuSec3OdleJ0U9DsMPvNr/0JHOOtrmIW3tkJXLfNjXFe4Gk/g4zWcWWpp/xi7he+sJ/O67FdDaM
QCuAnwYHta7/KzNz+eNsqbXchnb9txvkdoX8r6wKc7Q3qaiPj6JECzGCvLmP8Twf0DHFARqEAPMY
lT5L0DKAGkqd6eR4OnMKTaox1W9IQtcMaXyC8myiTueZoQxXF12fNTT1K921+08/RhSB2pTou55l
irqzRLzRxw5w3Znw2xy1w3aA9Oi1m6oMYBXt3zDSW2zzomRJ1yc3uljQRYIj6/B6bhOMQ2cwvLnr
f3T0FIPG3/95jtTXtpqBI9KJDcN5JEm24I7cBOEL/gK8VlHYXIzYOqyuwDJTjQojK4gXIkOruuaL
tttTHjuRCAlltb6iZf1sFaEUXTAyB172xY5wcpFfMjW8l0Vx3RR6mXHbWv1TNcapcmUnzSKHkQ2F
1FkJerWbP9KxRUXJikV+mWSTzVL0ngEj4jMvDBpCfdRkuOnARzPsXXRYWucBM47MVwfFkbR+37Rg
NuNgVyMBRY6SJJfteZtLcFo47+gxeh7bVnpZuInQYJ7GityeoPNxrVl8NflrLd+K5d9Kx8/YaPHd
Qmj0DZRqUf/2PczQ9UtrM1rTJuDhAVssCfgDh9KK/uqay1Y0TVqAkiIZx8LLbjAZTNBhhz3iRhU7
R822X1zTDQxf1zkD5b/4mTnILbQijPlSqIJtFmCQRw4yya9CjuEZ1I85GanBAq/wdXSsfPLUkjIk
5+EbsuQZBiUC21mf86h72tpUG316pzOiEhFd4ckez22Qogky8GQPiYTOUbqp6Cmby9zi1+luVWAk
a3JTOLYvkAxCkAgjGP1nAx+xSLqn29Pyk2oQcWSFb4Z9jEvDeEZEUqu1EdGiAGBLnb0T9MJ3ERsh
skfOC3Brrd6t2nETnuguT5lN9aakLTVElzjJZyhyv4VciYPiWZS70bpgM73GKlzlSm223G49V1yx
H8RanXKa7WTFMch1AzHteklVckGgOyzdUe/tECM2lznu7kVsjza4o19hAd43qwuewMdTeDoFphqH
4/1noBg1S9Twf1GC27tVwsZENvPxRgJnYfWkDc2XiAHJTqDg7tWyhGZLDOobIvGHRDhQCqP4tjlW
vQU6nlVLIscji1WaWG5EPWYbdaF6eqIO3z6ZSw6J8Ox+JAv59PpgMOu9Pe5EHegmTjz+IhBwVX5Q
Sq66NoUyzWH2+JuL0vsh0aLnm7r8GJAVarkrqQ+n4sE03uOWhfqH/TzWujnybCHhEzdka15wkpKz
0c8Y7JvgMfC5y6hS4w+DGymqEtFf8z95uziDrXoRRBUZf6DwGQufl2adAxjNxhY8wnLB42s9Qgc0
Mf97idPJ9dNqZ4da9h1KbLgRYtyDQeZPETPtRcd/xEzyEMRc3WD/5fD/MjiUkTVXoDiLbwT2N9jz
PikLY+4JTvrbIY4INKdGMMTVh9/cji4YR6hHEewa7y5Y1gFvmnbcOVngTdWdSSwcRrWkRldbS7De
Q0FggP0ow9qJmJ4w8+K9O70MFyC2qDsetHZB+ZKyyVP5Imd5+Xrlo9qRQ7vpqxUJupcD1N7wK1Oj
U4mfp3gMdEE6zsQ3+g/xdHu1xEYAFS/vQtLDOsLyYEHv8kPitoRozWrEVCMzbC8E3DnuwcWAawMO
bDupYGqPuq8zfT6jOA4/9zxU/QpRU4RBCzi8nzu2byD9YFLC/Dw23XrZrl0CWOOii+DMqoJzrxOq
iAaQAmgt1zmeF26H3cPso5Rb2Ypwsv4e63c/9lFuN1lxupkv8Mpxrt4PJ1KBp81NcOnhaUe9vh6M
FtWyu+ojrKjD9YGqXU6s6xPi5JD2RwTSNvAPms2NbBOkFEZp9NdTyi/rCr/2egrGsMHjb5hRPR10
fZS7KXMs24HZyRuUiJIeTZNAitP3MuzK+WAYzkNUfmbgYJ8vrutQoxR9A3B7WY717po1ss3AvCBB
i6o8DXqW5H+VHy1bpDZBQsGh6r6k5vfcrqfMwZsJZluHq+oxyHMHdlTMu6CX0osonR6Ix9DJmFyK
Ja09K+5y8gMazvqCLaW/1UicStqN/gs6yjOg7n8JbOGcuFoWQOrgCK00sxMUHegj538iI1sKNeFT
/PGd9Qg1OBu+pKAXdb2qJC4hsSrVpLqMilxtnTAzTu4qQ7M3l3fdkAiJXhz0zQm1FuyUD43C5P2y
OYm5RJBYf3vj3RQJKbGBdbUFOLdCKH9en3q2kZIRnYZ6zCJxItuOWRYnB6XyBbWStjAm3D7ikt4E
UX3WzU+aryssjgz34hEsiqIWgo9DI48FI+nGu1ZAaVS9fRecFrUN35n+qqC1lVTTnEWJbDWLMd4h
vDTW/SmQTBBY2jFgP9Ayl8NrnMy4/fyMfdkQdir5JmhoCdCwuNn2MnHdj0b4VjjelA+jY/+YCci+
HV+Om7iEiIhk+7VXJ/BvTT322uaV6dEryAfvAasVDAHtMf8IWmf4GJSzDK+iVRuoIavMLB+jF+KB
IpSOdD3U9Vab7WPUyvLiG6WiRDW91CK+G05TU3IP1c6ji7Mf3CHCKPA5Ib0fzSLwKcgqs6EAx2cT
dgsmyWkLZ3fAyjHfV3XkeqHzWbkhpSGLFOidecUv55rw6ET+20gE3Ri0qLqzrvy8UC3UvnKAMZe+
ZagV31tFwpdFek3xbOPJh14q3zmQvam6VD+UaoBlkaUOMQK0QZDy1dAamVm9HJ2Mc9m3DMeEPOdC
V4QWN9esPeFNY6sw56RDlXDCOH3z3jZEcKSf+eqRFUofB3kRgx4CcX7KWKJamza9aT865mbscnbl
UH612JPhSj+2bmEcG4ye4m1IxRKLech/JARt80mywpfpOX5g7S6HslRujjgHTWQwCfGflMjYFcS2
bJxXwVShTeWybulVRekIQgvUvTBPR849KTQ/FIaCx5a6RVHDjf3VRnLYfzm5F1dFvyX7+vSfoKfS
cDIHHPku4glnPe2AFgdA/CIhilVsdwnK8PL1JBvXSDCFZ8d9RongaKx/g82RhBjMnu/RXKLOYZ/b
j+nP5p1F6n6Mkk5mqWljLR1RtvaHugSW6hiP/SF/s5HrlsY73iPuT1jkE3SXn562v3d1dvwxXd5B
nD/RdFjfWC0/HjtgVBgrC2hyT0aSzPErIEQbAFrYNDMYicqLwJOqTkjjAgKaBqVFTBpUqa2FHJpV
Uow0djqAWYS2nLIdsJLjaHNyvejn4RzeB2XivpwMcPHFMCui15zgnXase3HiIBR/5moJr1k/6dXQ
jAiGkaegswdT9i7uWaloFbMAZ73BvDWTu//CNL5569PM1pzH+ZtyWu1VJj1Bwz5874opNOxvyehd
D+z+E3E6dcSrj7GuDi2N2TNFLwq92C7l29r3+/YYLBlWQFxIA40m6OhO+KivZt6lk0cWTIRI+gHy
DH0Jfn5pvVEQ9DGGL3vyWYaZ1avczSBks3z9y60hFXVo9HyFjP2M29x65ME+kXDiximeOqhuw8+0
oYNAluTPh2HtnuF7W/TJduBN4RSRwXjhm5ODdK+lBTotvMCysIrHwGaWStMDk1OLFrhnY3wmDLuJ
r+OKfMJEPy8b7OBeGsfB3zmxE7W4/kj2rPjf9UnPzGXMf7XYc5hD2Z4iEkhNxDTpfM08PxCFbHlO
Lu7pJSCMx7g/1gABUCWhcVY2wHF2dArfmL3aMcKbzkbH0rRoFFM11+Zn2ofWpF0dgO7YqaTog6VM
cbEku2IyTz+6wk+HfPKGUpXp9MUXr9RFy6Eq/AcgYYmrYkEYZhUiKKspGpE5JVQeC8BmcuHI3O8t
DoikRbqXUuwBTjygXPqcV63zO4NKURA0YecMRrJgkUiSSWJpF1okd0vAMZkenSnBWCFSCrmk0AwC
zr1U+I0Pa634k+1IQFF8Jn8VYWv6FZeseCJQnxcYU5qcER+2I4BmwSAkjWdaxSvwK1UxXg/bfT6k
kBqvy0e6W/9V3swaZyKB9EzavWylWak8AAhsA2w5dPguWVbfMFKQ8+Tp1Mb9Ad6EDdTNiWnfz6pr
JjqIE62aatD+LhZIg50NKWF653efo73WGXPcK69i9OhYDsy2Q8vA4HF8FlX0p3RLwa1MRnqU8pdA
xxUhTaOS6y2f3EbcY3OXh/gLTng+dwYc4cXeI5Iw9fb2QOFY2UXR9WmIuNLm8YTSUrIiqmZiV8Dg
AloLg9uZEgFuxG0ZgczMhG5hxruiCYOGhkSZ+h56mjdy7SPDGetlKZKrNmt/Qirzcu9jUCZ2NMyZ
/BT9A1ORow9fyIS8aq8UnxfXOgygDKCEpWNncsmamapHQzNI2ysKEyrDQZL2o9prrYFkUURRPU80
M9dypMCE9kQHAl04CSi6Y5r5oAwH8GKnuHYuSkgb6yLRW7Ga9W+7jUqZoBtn+MY9C8JkiQTiFeZr
lKh7ms3LQr+U2uLhClZy6MIPlbll+41FPjpRa+ZY3AJsh/9yc2yxj4zlNBS1XGwlJQktZMVKG9bE
qbgVFOhdXBN5WoOOYjWd77GbbW31QNyzluBs3RpGrBC28FldIxBQQLuzH+/4AJwWmV+vNcA6y6/w
LU/zMoWWSCc8hiHygk9/JUvY2fyURahxbYOkoPZLYS70c1EoYD4xiH8HQq+4kOV9RJfYC+LdVwom
Rc07JMaBywi2BQPAXN6EG+3GqXcTGjdy0XeiVudihDxgud6Nrjvuj3Y08YWKjve8lCmwseXBI2nI
tlDY7SBqvt6AF6w8FQO68cGLuw93/mhLbU5C11XYKHvgKw++oHBTrWTGEGn30/YZHKuCBMyAry9d
aD4/IfMoLfAQs3TqT4Fkan74KYAP8Vx3n442PmqEgKBLG0wX7XZjQnFQQgJ621Al5MC5WlGOvCVc
WQmUehXorr4dAzzqwvGbBwNQUpqC6e0PXcF191QKXIpRQgyr9f3PFT9sauXAtirm83wpRCR6D163
w2x6D0twHstP41/W+EDhd1J2amLoMh+Y/uqPA5NJLWOeMZQzwWBe8cv2LZ2A7DWFHoPd9cFxOBCD
7luklrHk2ik3I7As7Ofji0M6Zx8wwhd9ap77MhF4qEbDjeVSOCV2OXvhgdmE+NKWApP8LlETEgJn
FwcF1xnGeekg86k3qI9OT+ZKDe7UrRbnrncE9LSkGozSJ+uZT3JTDVaJ2DyCi9iwHykr5/ClO+eu
y44doq3vOSYuddSx4j/vWdvg8FQ/Bk6JF7aDr3aAaIHuIHpxESD6s7/sYLenkwgQwLqS9nWj8cs+
4OLG8M4nGHCF21n46jQOba/U4z84dfIzhEpPouLpWJB05/vY2MRQicic9LgiHnxqS2GTPzTaTs4n
G4Gx0a/Cd5VTQzc1Gsgxy9M0psbUjB+eB6D3dUKTIuJldP7+3BbM4XWR+U97houKreLBS/taqLmd
hp2QL4t2GTvZAosG2o4DdTAi4CdVXfkoYkIEWFQizy6cYZ7UCOMcqYHcXNlvLoRo8traVTejeWkx
u6TfEI5xzAXu3CAcAfP0nyXC1ry9uh0KUmb5xeN/nuUzvN+0kgbDk4TJzUeRn+JPExy1XudxSYgw
qba3z5X65l24Z1T9pMLbKNcyHNq82sVmNS0wyrdpuV/IYhKh2gkmMQIgrmJpD+pMInVj6+i5Wnsy
LWjv33wP6In7b1TAYkZQsXQ8P7MXB2RNcv6CZGd3jxLZoC+HulPoALgAtY7OzrLN5m/kd/NWuRz5
7OHuQ7d5h7354W1chP9S/h2NBCBCcZvrcIf9XAhTBjHxaVzWezzj/Ux9mRFxlvLbNeUpusK93rLe
0UY9ColoDe0jeUjM+szAwA1HvJgn0z2pigAbbLWipIxB6X4f22VpkgZNWZvUmXud6PULTx6T6v9D
PI+yTxz0NisUGMGXM4XeyhOg5V8IPdvdZEJY9bLhHUPycFlwTPKVE87tYJhn4p5ewQKKiDEmPYqq
wK+Y2Mbzx27RveBHJl3Ap+G5Hf1W/NDu4bI2DgtFfzO9poKxIFZ6GGJLQ9UU1Nf9iHCzWN34XwaP
MVziX2S4EQHaOhM5n+ljrtZNKr9XG+Qr63eyX/kMO/Hzjwx4aWmG7J3O/u39H/NqqdHrv1rIvMTC
Vu286+i2+X3CitNBM/xjKTsJVrLp+QxDVLTzqLyS291JbrzBeStRuG8JZVYtrouZE0q8hXdti4AN
e88l6oTP4pBD3mHP/fDh0FLbCT30Ax4IPMWJLoWvyfiPQLnGHLRXMZtyAhVHaIevsQRzRRLWfUXA
FgB/9CNyYvYFXfFo49VZwvX+7OfYqNXCfpWVoySxVS7F8aAMBiZ61bRUXa6HCs/0uJF03+5E/Bq/
Pgyk3jNKVoZzG3tj4o2yu4xD1nmF8+zjIUJHMGRfvt6L+q0VfEXXSPh/7ob9KGQvVhi559U9NxQs
k6OzP6Wt4bS9Xo2ZFDxDbjrpc2TK+tTRhjrLXvCHT0KGiZgKe+ITjecHHBApqZ3Ed6dKLxD6M34u
3JqbQepy+tRMkmewo9Cv0gTB0juVDSfUTe8MHs6KfEa22akM43uwlnA7V2tZ0WlYTlMohtCfIYH9
h7jcNNv/FD7Ks9L99iLAy57+RXO7LoFdNXmCwpHRo1c3/QuHmIekSFJbN4+zudR+mCWp7fk8+kfK
oYFOS+exsD/bfx2Jrh8PcQtXYfPRn45jJTtTi0BrQjZr01DFVyPhKoMOieD7N1wVk7IyrZPDKzIE
EQoSLGTLGQrDllVdpujWfL3ztohYxpbVjhmXiNoVI1Ft8sx+cu6dlb5+t/AUK6gC1dO1IFT/X9T0
vJVpEFdarZzBu/eYhmZ7Xzy0EBnl3V0Iw65oSHayK1WJe1BX1Cc7mX3aDrjVaYIMg1OSqTlcWhJk
lSORc8jj4KeKMe9g5Z0BLb+qq1Sfao6Fub9WIr3ZOKa0uU13n/ZphGANR4pB2igtoYebN+A/8mrJ
ZWOEDIOFWCC4lD8l46d+879xpAwooQvA9P3xOzciuRs4APfyYL5d/HUR+8SI/5T4s4i7ebK72MTu
nmMrEdPiV+Om2eWe+6K8nS5/II2iR4zDGN0NvQfke4kc+CN+ufzFrw4VUybakKFwHHFBdDNVVB4y
7lWCbcVRIZFS6UJB2mL0JNIqLp4F6jC7s58a48ssBy3UobZRj/mFNNwBM4WjrXgn0R3OdmHmEw5H
/+tWOfugzWRWJlKsVD2G3jDwI6TXxbS7gnrj8q6SG3qQseNuqk/3KUM4L5qhOumEvqTL7RRy4XEK
QwlNU7K6Ma4Mq87lqErHpHf2FSPtVTR9/Qjyiz/PNx2lYBgmim3upyJMC+HSZ6+QAOIwNnT+m9F7
BTtXE9xj6eLpg8QBiaLU9VGcDmaiFsNiPXr5IH1iE0XkXn0h2FaesL+G/fmsSbfUit0ZD5p/YyHP
lFy5uaGemN9SMq1JCmi5Wriek58hQFl9TffGG/SKZWpsvUVRvZSU4rDb/6pBevT6HxO/o8bgZonK
pKntAKWbiSQhMoqTUU8ugfzZfOHKpg2wauNOF0bmodx9Uabxl2S+NQKPvmJs2L6Md2jj+iGYi4vF
AGLCv/63sj81HSilKdberoRHh5jbpBRe1/+u4+srTbBJjy8QYf5Ib2STK7BdNoPjoXxGpHp/WMO5
AP3tGY6p1Vs3/wqVlpfSjI/HHq/LlZzPSTJMYhe2dW//nDeddOi6XKH4okZezdYxHL0ERqpDd06G
ZFP0LwdtfZrMNfUm0YQNVvpc/qgMGIHZNPdNkCNzSMQVWy5EMomaZKLGX2Ii+F5Xf9DitzGkcAW2
x3w8RLTjkNh0Cwd4cBPGU06xjPxVVkHOavkSQ+HWetwJw6RfVPYfqmeF3BIrGaaHbdfoVlUJpQuA
0yGr7UCNPhucc1oR4dJgy7b3ahwE8MPa6N02vMfuytir2U6EJ45EiZ3TlyAihOQujJ7AXBPmzVoi
3P0wdwxa0fy2VLUcHEnbQ1XQO0gz5Cp67QkByHNi4zfUnRpyreQraxOqO5DMvKvtJ43ogsRBWhaX
bVoQ0XeYHlf76yaTE0O9RE5hv33hX0op7zfRoTcnPa0FeISyntjeKhJcsP9pWQsCe9+xsLG7vqFW
K13EBKVAx1F8ACGIuYLd2n0GMvWwCSYn7epRIelYOZ8w7HpPe2KWX50rd128JFjIY87FgLqWeTxp
+hN0MKTcv6xGojJ2U+8TUJK1T9YvH+Xvz2fKlEBQMMkJSOohw/jNzOwfT+nPAccpfQxCfdpQ/LD2
i8Jb+TwONtS9eNLJphSZcvDYW+raRLBKYVupbj6v/r22umdMIQ9vSc56VK6IbRImnqfEjHtNwSkw
PM0NHhA/4uSxhKBV4M4Q/VaWnqcwkJ/nOVdtBXgFy794ipRJXG41Oep4yk0WRwZONW5bhZIE9keW
taH+R2C/gbv8seNJrwpT2BbxTEV69a2cDzxPHvLTjQKQC518DgwZSOhigqqLdF3InEUuyNj/X/0Q
B3wt3Ke3YTvooOez/7M1MT3MhOCy7a9JRWxoqPsB4fXs3OFQ9NfnkuHiD/N6CHevtp5FxcuFIuYj
l8k6AXZmiuDB2LIDaKAb8lk7PXwV+P6zF/VfklUruP3hDKZJ97wyhlKdS4SUC1Q1kRvlbm5xZRhO
sXY/YmLUpLZBhgct4RC7CZdZ5LmkXOA58Qo9VTPDKg3oDOJtWjX7QaIn89seR8TOoXxlnrT/CzHZ
qdPTYKBNQF5ftEOqreG/vS379njKNA20j8yrLPMwJ7uyXkOWigPOIPTqfKf/asXSx8i47fFFUHhd
CHEVXD/bzlc9BPjCD/mrGlUC+0d2yHkQzLy6Y8GVbkZJ+xXwuxE+nbLjkImAO1Kdk4KDAVuqtI+D
MQSoSCwdzEURA9/L10Gf94DEDleM6glCX685JWX9rmRqFPNZlukMNV6c7gVo8i9kDYK13UBtNGR3
8RHb18QmHH+wzmlntLrQLqpr9bddvT15JJnMoJcUfn5W4COBSU1RQbXcc90E2MvqUA8WMIS/ik7p
MWlyGeBPkE6J1kTqzhiBbRSLMUtjQeHk3XX6E9N3ILpu+EhcKyMQjQqMtjuKKozmyWuSL/Tz4TKl
Vy1ke3Ib4f/E0d7gA9xZgplzWKlyrSQvkx4yoHC5lxVnVs5VsM28PUe1TQX1uVtCI0+g1wvd9dAq
r6nxylsp0ffVJ2B6GuMzSkQ+8gMUFbJ3/rzef11OuQMxNRW51qs+vz3pquUFauxwYvskgKsUW9G9
BJg352sKCtw1xRsBcANOlSKk1ioqlYuFKhLt862BMn4w7mHJDbP3kbbwylECPQ1nW4QZ4kvcZPnR
od5Da59uiO1UOh/EbPTIBdI7YsZAH6e5ikIoXpbu+wPBSs0+T46zCN1chcFkQUqxP9nLbmmKkTDk
LCYyW4z/9t63+v3n0U0tRiSDcSBsCUKj0Usrr5UYR63ZUQ/0njuq2PtgIW2/LMW7fz26E+r9kKum
Ai6N8WOIIjHBG3mkt/fjJ6ND64MtE4EwbhkfCAOWJroeAoPAPvjLGSVfrdphsxARBVFDDbmbJk1u
OX0K5lEBWRMR2jl72Ux6qjGjL44W2Cq5KOc9hD7anU56OS+zQt2ULamH1KpCRrn3UoJooNjcl0/r
A2qYSMk6gpHbDyT5bSwVhbtmDCiW+co26NFLYmTAYwgjBPw/Ywiv3k5kTuAKGU1Ty0xLyXJZcv6Z
3WQi3O5uo86rpA/x0O2uGid9HAJT+hpG+2UAGj4lK1VW1GHkl9rubpt5HIt84thcohd2YSmE854H
sWj26oQiTEuXTT5fzJURAlsH5q2JB3EKdaevYZTawsYoM2IOrajONG2edk+HtKwAyl6+kOeDj7rQ
0ShKUwMyjwX8IioTtYkvyVOM2/JA5xMyOrI1Rx+CnN+bzTsgDmcitWlWpihnQ2VQu9XeELSgkhLR
McvNLYLY/D8N6z8SVZt/XTcINDNwQRQ/V6LJB7TsASynww+4W61T5DxKsVGON/e9WVH7J1RNv/zg
gu6LKapE2aYsSjbXUpHwpcJLiGBPnttrfm3F7IEvAB62iF2Wj+9h030r13pSZMxXn5GzWUruPRiq
7Rqn+KGGHp9Cpzo00/R9lDnApLs4NmYyWdUeYJE7nyYZfGO5CXvT8F6HuI2QkL4kB9MM7rk1/QvC
i3J0l4LBCa2nPJLm+7Vfddtt0nvU8/UA6JEfFwW7kJmuuZHKy0jrqJ5cOqT7n7q0uFm43diiYIQa
01trfUOnoMCDISYjwu3sgPaPhUys97MHSmecFSF4gwzy8jqCLkD7uqGbPC9q9PMKZ/rmVUUu5YXC
HUIS3dg4tnheqLeOxRkumgskA98QR1JbkBfXXWn2rirciudlByh+5FBMna55RhGxz+YCIo7fDmPh
G99KTIb2z3ubYYKldw6gr3STVMs8AYb3yy9l83DOEYLltAONJCyA9Y92VvMjRR7BizDyxRhk2gRZ
gx5d8JxwWS4D03op0liyMSuNgIwKRmPo5A/twX58Hhetu6RGWq3ZEC6VEy9Ju/abISbHBUpKS0ro
7pvQbY/Rdjx4f9Zy3f3KuyaFhi7i5bx6RbCu388ioJv7oHmkoa9YZmT3M+AVEmgs36eF9ti0H11n
p39qB6jCKtXjOGdLzTy19j6c/3s5I68XZGKuzTeY9pObzJvo1xV7IJ151dVHm+C6/c5cX0GSZnxZ
IT5VOrLERmlOLSwDD2hRflWzQuvbG7bblPSB30CWAPpS+OwrrlK1hyqjxL0fTlzYl3VfIOIZiY1W
Kk3SnnDEmLpzd6v6EYmH80cq61MWSZhn/jn7qJmRqDUGQlCBnJ9ql/J/XI6RNfHgg3tZ+FWFooIe
dG+GDVe/jy8RT7r/89Hwjrc7BVSN7BLQoH+OpjDZfxSxOt5yfLjNVhf03dIjvsks9h5Gl7s7ot0g
5P56i79o9ar04BqvdFdPD9i0f7JgeQV7na1YmWu9+wkvgolJDdKC8qX0pksLSgAuc3E9we1hJ5O1
CABG2epJ5ADYNVB9WZeShRZ+CMpy30H6x9LHGUyqwKHlpKztY0W527IIMK8vhvbyPujObbhluFx8
fIqWzc0mFvORsvvafXnluIZ65Dj9AdrhPmWD7uWzl7dWOG5C8nmJp2rPOCBtJbnGLjiyosE54zcH
XGSbEwSMR11OG5RLKSaD1dEN5ZSl3Es+imZyf/3Oxr3pVWC8c7FwpDhqsVudBi/1OnYODaMqnSsg
KrrW8HsizGH11D83rIEVWE1OoFjiNbzgtW4HisbTAzA1XJJvsYo1FMDnZYyiEyqbDerELbekHayw
mcysykYd/1HEAhat2kFqhSVsRumleHsyNEa8V7/EMxSCguPQAKpObIXCUsXHY2k2meGXZUM81xdG
uovO/0zdIZ9fbsXs/wZzXwhvySYNId9chHqL3sINK26vr0vMZnIhy7iI8aEHkdSplDYn+nZHH46q
B4p0NimSJyrQb905j8ioQcf7fdTMY/ogiBFwDlo78AS5e3JB9dqqAdllJRSIrCfZiAwXuW4+94hk
seymwlGpNpSf//CW54F9pP5bi4+E3pmp8qnf0Gn7FOATVi6D9O1/ukMGywkJ9/RIktcOOUBquQJM
VJj96FSDte9oRAF9Eh+EunW4J1nZ/xzTZoxx5vqMnJLXpSE305tP/15+6SrjWAP2YSOllPKOLuMK
ixXeD4obyRwwnk4F/CP2gRRU+t2cSDFLiEfpzLFmvTKX7mTjFoUfO7T7OMAv0cpTl3209qWdXQ3H
bvXRNiu5gDBJigMfDS2+XCBdQRumdfE5UTfiI8YKxmzkll3GHf/CoOoCyzvdLNYiSDoQPOI246jy
T3tEqIS19+0RA9Y5N3sOYG0GQ/HtWAm/JzZqtOX1KboWiT9KYwbOHNpzQQssail6uLZwzco199Se
rGCUz0l74xCnPGecwmSb0ZfYO8rUyir/bNV0c+li3q4gQyiwanqEQLOqEFxZRPb+uadhdlRLT1VX
ARu96XE8k65i1yshYtDSJKKRFKM08/ekn3igFA9KUGZbHbo5u/7ufy4P7Jt053DTeCakH3JUKASu
WJV7DgHadM6ycLmnCCHtOLOS7OXL6Q7wLfs/aAmTF1XGl9q/+GPHjt2oHD71GFjkQOFFYfiMhNmK
f+Kw1szyh4OMQY2asj5S+V0H3i2jg1CyI3WanI+5Vp6IQgLGbCz83mcMcq0nz+04Y1BZBadY4Exs
iiZs5TjBJZoCHq2JQjUFuNnZHZKruQtLuNrkwivPqQteLyN5KL2agtXDOnOAT9xCt0evQpZkV4J+
Kvnf86TkyU+fKv7ETAXnWOWxKn8QETrnTk8FESyQGeM44IOleBjw1VdIFhcbzrWlXwZbzX0wUva8
kekeC65U4X9+8nNOHDQqf+LyR3FrpQCw1xOg60/sXOiqS1cvGMnGh+4fhz/Zuo8Tcq2sTrVHTb83
qEMBGHIPvajy6Xi2jHCwr1buN3ec2OSDCqC0t+a5XtqoUuGJaCVeoEwGbrSGamb1l/4rpRQsBKb1
FCxPjzLnZo6krAQtmMUDSDqPbFALGDZ7LG42Pu5rgSiYNLb/VgN6wWogv4DAUXC4ouRUMOUBToa4
xt+dyd/3JuCZD7JJNCuom5OyrisK89UmsrXWJA/K6Z3y7dIBS5CrIDp9JZty3/1EQed2gXLgOHXt
MoycxZjMfgw83vwpUH6HEKD//YTAVxDOGNC9u7zT2/+qNVVU1PNsBAb1rpt9yCqndLRJ7eiqiWwJ
tFozw2wMFGwXcZVDnI6y4BF+o6XsruaTjRZlArfnZs63zsXuNyOjtyhjziMWfZhhAHyDaC6naDPB
9JyZeYel26cAxPKLA1Qj7tVsfx2r2h1OmUNOVnqR2MJc5+lHYEB4VER2jOKN2Dxfel4O/kjvLNNA
IYZtxEqRwfddXtPvN6+ATYNyyLonVU/xYaazWqeUIU7hhlAce4k4bpH4J0qzgNxKgKtTIBDywYMc
FO6IHFD7fYH8ePuj9b4bRxvTtnl7zNB4GACJg/7mruim9nAGzo3KUwLAkrn9SECMhr14QJ/3kfAB
SspLilMsjv84SYbAOd5U115Dr0qca8QVIXt9FSciGA2afxOMxXhaoS3jDLuMnNh+Bw2ye3A7xNx4
VLO233zMYPpfxdOY4iSicQafhPT+ExiBfYhz19f356J879Pz0grepwIMOinZQMyVcDQzDJ1DJQ6d
oe5vtB8fvUWzKeyLB6nHDterIs7JKCsyFn26OR6Y6wcALSQ/30jTiw4/P2kOghLe96kri22F+Sxz
NBu5CsLOSvBgrU0PNgsBuGDw/KzpBa10Zk53pzfA68AIbfIEWu2KMY+uZVUEpDPJAdWqDXBPB+Tj
i9gXdDEAVQ61+Fim2zvFAdVwgaJAoEwXN8ogF8pkaWkCEaiKu8HlxgCYxnA5rxk41d73E0hpQD0H
afdAplaJyfDUEcUHS9VTUhU/L/XR9XTqdaRdRqTgw0M7p4ax2TEOP8QhaCzJ8Yi2VyR+sOdeJLXV
su1AgkErwoYmcXh/hZ8SAA48Xk4IaiOZwmmGGVD3hoOoqYvdjvmN6zCsxSNDMjClPk/k2JJTHPrT
FhIr2BW3QSInWPvl9372neNE4DDZJtNR6PY4qigE9B1fwsk/bQcjWvvs2Lp3XboB6ZCQOsfL1Ixe
I95qrTWaVHl/pylgcHULuxoWf871cIWbazLzzVVrJIZeS3y7ZjmdRRVcNRiwXJioSgLayEWGTBXr
3bJPtEJe8yFXej6UJ+BbzOQvCjCxghKv3op2IJqWxb4D3LPYUfIuIm33GDdkKWI5L3mp88nsqClQ
9gAnSJ2jrytNEOwjdVqB1A2a9fZushBm5hs4Ql/mTlh44JmwVvA7O2NZJEV7BXzxceJ8w725Ncgw
JspuVChkHcSBR0PcoPFA4yYi3SpF7JCmVq6ewK3vxw0NgNdU9B8fEcoLV0WIMxTN3/ny8urIsHAc
himJ7lzihqFJjlG3gdWcbXPhf6gqmuF58RSW5RBgKnp6Kxmw16zBRZaStAxQc+GM8tdBT84KD/GV
R7vsGXjBK9Y3yUaol66X2uP/mmz2yEXbJ86cZsOo7/HY1RnXwipRoGWqUPy0J/VhFl4Yuem9IbG2
qMGQxyvPoiSSlPxd6z3IJwKHHxjb9YFR1tClvkCa8kR8YJv2lc4ot24vzQDBEktbEddwHCRSxtb6
11pnyl3yxHqbKElIvL0ueZU+C42QKelX9t0ldPyxGa7cUxl4tm9uv9yYn3pnZ9SHa3pIonFhgPgd
u9UupXZrgQ3clRLnOt/EQVX80DnnE09Q6LDU+B4WLJoQaI0TNozQnyTr2kWNrwZlJZonkvP3SOf4
1+Lk2EJlqh28p+7yFwrSvRVVvzTelq+5FCf3owCL3H887Sh0xJgwnZyVzhp3JApFlLJBmL7ltYXP
HIgkDSMs0KFaMMckenZal319lu2i50S0GyPMXvSuOOLKj/sLbHHTQeUXXaIPDpII3FSGoKnTIEdY
Jb/L+luy/cg3ynoCfLQhTz/Nsvb0x0ruoyacM7Wi0Qxlt+CHWz3CGpf/PZ5+Q50MxvF0qNvcy5Kd
UTPZTTLnoFwg+HauKZYOfYsKCqzINGz8H/YZDigXZ9OrRO9MNEktQbmZbWwy4j4QcKvulxWYRppb
hUgbB+f0tQUTKy4JV8Sh/S8fcF4UALJwiNZKJaiuwJYJawqnv2HHdoxAZlUhkRS7qk373azFp57n
qR81nUMyqab3OruoH6wmgue/xLLSsnGWyASWXOWu9BkqzJh3kZwT/wNB18kOL5zF77kHVQuxmNBx
P/ds4YKnQVfyAANm9fSjciFuDQoFZYg3kaL77uVlBCxlSdDcIefbNJHE6VPwNRsbV7c9Q4lTIibd
kMZoFnt1AyPB2mBPlL8NkdJS4WqpVUV+FkJ6+s/vBxVXExHPmgGhd5kS3Kr7pI3LvsxNgZRE/xvg
wMkZiduF3ZogXsXKyibr9YfrtcA4u7S7uieP120MEDLink7eCHcj+LwTJPRJRgPxJdQg1iFWSIJm
nWkCMcR6anto0bXo+GDtV5CR1HPI5dDL2rumTUpBYrQoignfxguZc3QWvyAeTrfDTaw2g/83a5V8
6n5NiGfbUzY5WDbwn4hNtfOKO4QtUUuZBIEkKu7iEsIPl2WSq6DwFUV03Q5jF/Uq0aBSzZNovk0d
DEk3rWYLyb7yVsZjcSfydLX2lCht+PT+XtjLGUVkLT1ZvLZ21+4zFYq4eeNqNUIRlyMaPkj0E6AU
Uw9+rso6+DQMK2GcmWSX83S/JpkyYvUd0P3baLexbbGR4nOks7W+TiXgvaNlCyDqTWtIra55fzjO
t3gkuauOl7Q7d3mZ8lvbExI8lbuYH/NzCsfOhD78HvaIp7VTa2cYF5Wa3mWRqj66LpbVQNbc7vIg
5SQtJnFtDX89MX0qBn692v7n3DVakPdyprkwaQ8LJ7TMwSy93x6SPQpIQmiE4RsTE+pbHDQFI9GI
EXINRF1+uSw93tRRlhtleP/gQmq6dWRtx8S3QnHyCfc7JpYDjpaeYX31OBS0i+t93BXMzJdynkqk
tmgT81JnR/oy/uKVVr5r7vPmo94+1DzhPmLriqhC1sMbJbtdGwdyJKUJJcySZvy4WXyYf1EC50pl
8ANczKr/rW/OzuXsaRQ9ZBEHQ7j4wVCjVoMXJP4eB65AUUl+AcyTwALbvs/xP72qUNBZ57bskNrs
zpAJI08TkgTudH2P7i4fA3adO254wtOsWMo4dYgc0xpkUC/ZPwVfrkETAJGpHHdDTv7abuj/0pJp
DxB1Wge4qO2HlXPK6Fqhv1QAI43BO7dugXeHLYyzlOFcvH5SDvbflVYoFlwn9ynwXY1a4z2Yd6vU
mmwU3kFaq2tK8Mi88BzPvSclTpvOFwaIqfBHNkRN+NSg2vDy6UIq3smA9hnrcrb/Uc54IvnIUJ58
3jTLfHX129cNvQuIxmb5YJp+tymbCdm30mKliZsKetsVLitBavPJtUTr31Ze2ookuLCXr+VK898z
xXk+4hTlCpUUMHDXsp5qJdkSlkwWZh8OLzXFVLHdX23CmeMo8gSnklACJVkcIgdUILsDaLL9ff95
tRREIoHQtRuSYpfK2P/I98kQak6qcCsT72jd30CWdqBlwV1IPZatwwDU/+0ZoXQ08MwlozIk4aJD
PRTM0eY9y5MNwk++a9hZbJ6+rNXUgmS/YAgmwduhaYBjDuEBMEVLZLNdcJczhae3kOVh/pHd6GOx
3Z+SIEiYGjOO1a/3qZUEBlx3s6Klfp++9SbVSvxcqDEEpxqCDKGow2RJ78O90wIq8EP8mA1S9bA5
Nyza9dYzv218XoLUwSkANQFFjGTGQBT2WBrDC5s8mQed/GiMpx1edqXURPnyOQNJWKFAVnfm/qIS
QfQ4RX5xw7Kual+wzVJ7JqE2oHwrWiImzdHQhLjyF9ylf9Bdp5c6jL4A+GNKZVj8AyfpHDVnlT5Y
bw3hwLXjW1cY07LiwV2a1eSfboQedQpCrKAoTwioLltesGdqWa0YgFaHBW9ff/5YSZxI13gf/VUK
VIYp7/HHKKiXlTUP6MW9JzYNmQV+OwvTHIbFDLgtQv6xdZk/HyNNF4XGoTYPXoHRtaV0eI8mBwbm
sQ0fF0kqq/IySm3ZxI1dFu14UuxdHSgeyGHB+yuo683seVVCMTijrZ12dsHOJmDqyaYZjZ8Wjlv9
rahlETD0wYsw+OavVpVb0thFswzAbOryazp+5qTIhHEkvS/cwNhaSspP3KKUYlJl+hVHx22eWmad
reHgaP7uiGbCryURaMGTL/GB2AGAcrsuD5Z2FOlNLcKdwY2hMa/3iyJ6SedMY3f1PtqaoLSSDN/q
6RSlDp27VC15fjS6s4c/wwN25/N7dB+DJjlMDmXoENCNR12TTaGb8L1jZA+7O0N4g7B1nExyrRJ5
njCiqO+t5n//nF9xOGGziT8TKcINi3wN2y9BK0dpcp770jkxNgBbyJlPHXUZUeZNdJODax3wjimN
B9sCsbFvj/oGazVfAFS+drFDSMorz4s5f4vX026fgYqSNALUWO/DQpNmYrrQTSpMHDg682iDG4G3
9EYdrocfDZuC9P4rX6N0QIblgeb04O6YnV/94mMOR6tdAwVEAh/5lm0UY27rWZEqccQN3Xr7D0Ni
7HYIqhlY9MFvmeINC2zp12ONRubA2/AH72jNmrFPy0aXpBVpPTTSSYngEVSLTHSzy1ob0wf4F9th
ADjYCZ/9uIW0IQmgNTp6p9Bwbrox8m+Uun5QJZp7H3dqq2KLXFx9lRNXL2mRdil4EED9EkMYDC+0
hziMXGFX5HcGhrWKm43c2exVDrhNeEVSKODD+B/ZnZXzTGetpYTvYFeuwTwdPDkGeN6CJvDM2oyO
fCVNGlhdxPVFP1CVR0qQ7eSazeseDxN+EKjdO4NTjyud72IaqpLSMI5aZzzQnCt8jO2p6ar4bGTk
8tpPile6FF11cvN+s0NQLgrGoQe0HsK1ua354eb5h1winUMbtJIc7V19O9dfJRfwy5jD7/cvqqrn
pXwb7lvN7gjvO+5mezN9KEDuwvbcxTER4pDW0FHoCgxk1DaVjtcqBRd5iLE+U7BjWfmHOGlfM9fs
0GtgRXP9pTBwlpbEIEJAEIWJaSqnQY+3rF8BCMPP932PL9yBB4oe0K4siH+G0PdMNBZ/vyABcMrp
GSJeKU5vFXquxgAIMdlUHA1fWPcwaeW6Za0ytYnbg2lK3YGkkuSiFVGht457S9HNJgVgr/lWlpRT
Dm11XGSX6rnZkO3ngo6BSkzbKT4Sbe50cCe44Xjwf9SfErBUSdOhKOUpZd6+zELn4fv/f0m4IHHB
NZcU9HmlhF6Yuux+j0l0SO7VZBS0H7/wmYtvTdDNisIr7qSlbbusftt+qu0hw7vetiPgS92pzBsv
TBMLL79l6eHLz5T0egj/UNVI49HfAlrTMikU7a+LVid9ORkQY8ryoGgBhChbo80VKvUUSJ8n8wn5
yi8uZWnu5M3dRUDyEHUFqki2UwFA2gtWkz75rcJw2UThxMdJM3Xt6d0dPp/CwoFAlQnsCLjH+tcL
1jjLRNGFZGY3u6snTW/noUXvN3ZJu7qEJOZZARfkIX9rIX9B6EPhy3cKFooA3Enpmn02sQ2jvwX8
32Td5qiYwfCb+Kpy5DhZYam64zIlRH1w8TF2yOw+QsxlIKnUwM2ZKDnp9YTv8eQCen/rHopAg8ur
Yd+6vOuxPasXnWdD8WyMEyWH8R7kNhuOaw1Fm89hv6Dmoz7jxMRZnCRaagg0oWHvBrL7FX01Mrgr
07p7xqDDbBLAMiOjbSTJA/+mW2mKMKLJL8VLWBVjH6G0v6RAw6OZh0EvgawPUXw/tNf83HtfyaHR
YbZRVfXFDqX1RQMCC4oA+/vwcMoNeQ4Et2EbhjHu8nSpeEUJR7t6vGHIlauAqqjJV97Ix7Wo987Q
KjeN20+42bQ6bU+PUtp675G+25xCkZ0KQzpIelF05SHSi0p/7x0jQ5Qvx+ajQrI36pErMYz2viQ5
6lmIIDCcd+G629WxRHu209NPBkHqxWiLxdzbs3oDzIzhQz0uhuqGF5nmK+BEZHS46ohhdGCfQq32
lDa93kAk5aj+BlW4aRStXI8MuBjdRlnTDfvg7GbRfY0rsp48tTizRBY3g1nW/WWYLBvT6/50873l
HLZPmfdLtReueJ1G0jzAQsVV3j5GzQ9yz6OdXLz2rJNsi3fdT4F63uCNVkhG+6VQDdgrc0ZCc70i
qoEDewBUQhsKBAa5rm3elVvq9DaRO7PkAp7vZc6JJl/ZTs9M1t2r6oWHr05EunfRpE6ngYADLyBy
ctVaND6NE3ZamH/0Lwj+XN0LxNyxKBWd7n7Bru+PbFLKGXzdUb4wiwjzBNrBXyDeb42mI1YvZZLl
BiYKVfw4fhMGNBEShrUdNAgfd+ZDL+QoZQ6D0Ke5MgephgT6sOVoBJ5/xuuy+HZvq9DhuEW3X95b
plxd0hTS0hZnyExBKLed/dRd6pdG9AyTyIeGjviD+N6JfIdAGr/CMH85GLQO1MZbAk4VHcFZ2aun
SEK3+MZtc4qp+GiyCmPRvGGwTMo1cmd5ylzrMaU4sCTstETZ88G5my6peXoflmalAFnZ35biI2Ve
1RHs+bHyLfifp1XDmxkEsaICgmd3eROseluNcrx4ZCiAluR2cOpUJZFzwHMnOHkgy6aa2kyW/k6f
Otbl9NmcczhyjF+A1yWYDjt195eKZva3gHw6zqIeMF/JfUdVOOFv4h9MHmhwCyCurtTbpzOkrZt7
l6vKz4y/izko47/7mHOFlWIkjdZxDntMzzuOYZHKW9i2eJBN3RubomxxFk6cnmSpWEIB4heh/kzu
lT78HvqLKDt0eO7b6fjXv5yw/DK33xOdRyEizkfaXjMa9F0qO2SHWCrEEmpI2Cssp1Z4+io+ZxDs
FNNkUOWXi4Kl1nLVQsAXkFQqlAXDt3Q4mhlGuvzFFc3/xp6PjAdk0etgtnb2UEDejYFdhloNCHK+
UufeBDJ9wH1Lyr06ihZtjFe+skvV8XuMQkU5owFqcCWl63ve0rVdGQx7bzzkFPSBvWC3OrhdRKJg
YZZz7OgkkQt275mMfLD5eX4QWiM3UtfK3VXlIds2DvYaRUXYrxEbRpSJn/xxXq9T6hh++l6x3BnV
iPVYv43oc95bIppke1KzDhU3uXL9jkWNcu5A0dn9GtJTCtCu60zhzlDmO2oDvMCk1gJc6r3GQYlI
x4PO4mjoNi07LYg935nrdJxjzSnWsogn4CQKLk86eOdya1lvLT4YEA/a2AiNSOnd3WRYSFT3BCCa
hOhBMa0pLoTQy9qMgdwTDyfUzS9oO9dcPh3n6tsYI7vwhtN5fSeSZQRgJ1hXZJdq7oquwTmFlfft
JF6C3rtY96COsrs5ZPiFpXGJUdj8y8XeIq7EJDdPvwlFhWtGDuq+D3D919gtxZW/KWp9wUgMSVQS
1gTf8zJyGsMbLHwJBK5urn4h0uGdJ5oGMq8q/vwFvvAVjRnniOQ033x/EXz2KUdDSlLBhh0M0AmH
TS14cSDtsGXWx2NPgkbDPkT9cz6ssHyekAruhtKQlfyZXkOiS6/Cqwn4BANToZzx5vhyHu4mmOcF
yA3LX1e63qkpXUa1pHiQ/UAo3XQ5Nabg26zupZHuOoPKK9IgdUsM3vhHXrQdbzHhatns6jfm+w0p
+eOzDobbIg7la+SHY0Gta5LbqwsK3HSEiIJBzZh0gvtGYAxwKJef7VzQg5Yhtfm5I/1vSqx7fDu+
PQxzbZTgjUmUg1TYP76LUjDi6K8ug14jv21f8cyJNBh1Iwoi4ysCRBnY3v/oIjbZD9fVTZjp91Hw
wdh6zwdJPH1ZOuSdQIe/9vMuKzsHKzEwkkP/WPlh53lvOPr7VzzR+28HNPbq+Jwm3JMFw5UncmCz
mktwUHhjbXUQjsKH34MhynTqB+TICP3gxdEt38fyFlZw4NIHLIukj/KFsy0GDvcA2NppWhF/mmpH
njbrmwCJ6yb0wjHiGR9zOA+VmsFAVpqUm2zqorP/mF8JGACdCAj/27pNiP6RWXaKaGCaP4lXVSu/
z+kxXQAm0afAWJcIj90roepSMyTtPtVMixLQDDTHM8cRhuKcqeAqjzhB0GNf6PGgP8p9bKUXwObf
/C8TuhxfMI9X+NGC3MyzqM2insUcx+RynhhqSM+qj8xOctDfeGqhOhaam9Wf0a8lfJk4XAe86rzs
nsbH1Sjd4Keo9k6CBWVhvGbCb7Ef2XSGyhiL/igrJggcj2+DyVatJg7A3L/ykggZI3kA2znw3aC+
QO9z7aERoKDJZA41BDbMpWTOp0THcKwSVMwsKbV/zfe7NruBqrBjyWNy3UvETNMolR8Ej+GFV83s
ApCxugGERrrrgN5UnAwQQaXF62lHTsYSP8sm/pCcg6rK3LEK6gGcIeccKgRe/hMOi1orHbAGZOiC
eucWUk1piU+ouvlVFNGYvmzxNa+dHfEjvzCTw5I4D53jrhKlQY6EHKwoSxGFPxuxx2u4i0H6TIxG
Sb6RWi3KVZcwKYUEQISuVvTseIj+X6ILANTv6sbGaZT7733xigEClGhF1dn2cIA7pjPInHCTj9kv
zMuLV5fZ48xJCsKYdzQJVzYuf9rE3O2U320UBEjbc/eHHFaLGaA/LRPEcqbFgtbKrKMQQkFuA4Xl
Bdp7RMb/S5JACv7SzeOe2v1bsgYUK2QEbuNqM1Xvfcf9IL/HsINbSCkdRH5+tXUuV6YSiYgzrKmY
C6QB0JUpz2N/mJXaAKtaxAoH6XH8e8KknYyxeGKQOB6eQZv9puVtM6xzQ0C7aTO8h9vR0tcyY2e1
X3cyztC4Noox7J/2K1Kxpgk0p7bRom3g11Fqi70YjsarOpugsG3P1sjJbV0BFhZEtVPUiAMNq8in
wGP5iR9YSoITId2CM7fBr0rK6WRnxRjNUqW/gz+aWh1+wgEJYXefvPoE1pRjaT6s2WpORGDdT1+E
IyDa+J8k142JzGt3Im3Pck3mnF8K96BaxJy9rKNmpylvLuYl/1PgdUgucPUI0JfSM8Wk2QHeaokp
hGZCUo+aZCCA5+ZjhVKbbVwJwlNyHMohfqtsg16WccVHvEPNdGkzsdD3ZWU2zd9qHP95tDtvFSWp
mqP3O76qGVfObQdJpcv0TMlciJuDjPkuRn+iccYtbWhMcefFHeinwdorSLh4lqyumanIiYjsqZnA
et+kMbKiIE+tfcDu/LwwXi9cjv9dyCcrY4+YgV/NI935ypyRRndF2Ucn1+T4+5vrdAMiUd+QjOKl
gyAa6RCyI+PZgBMcnGEjqL9PcYmJZIapskFi0Hgagz8U/ohMmEaGv8ZEehVCWly+b0Fetm+jju3o
W2LqPg+3S9KBHhIpHYZuaTHdXau277YJtP5acv6eZ+FAT1CAJxhcZmGbwCZsX7tKZAX4kNJhPfhI
wMxHJg3sd1CahljudJDiZ2VoHd0KEFbStDKVzm9JbJ+3Jol7CZIUl1TNKUwz67cEGYd3vADjjcJM
KoMUDcPT8Uubs+YrLlth4toeq/983RCjJsCxloOBuE8Xnrfvu/aPVKu6qtEW/xqEecqhBQTizN7D
Ti8O7GdQQEvk7z0iXRPOjouc87DRjEgoFwRHLYrASkIGFz4Y2IiBD0Zg7CROGNXw0jchpXvxMAFJ
30xH1C4ZPK478xdkQwcAlYkKSQ1anuLbi+HRavpgI6LNi0v1RapGNyAaDOsxYQVqlL3dqDj1N6MC
+9VYU9GdXbuyBQqwm922YYhdt1Ym8ZC9Z0banChwB/gMfy0+A48I+mYVL8QCIGFxE31hxAcjXL0+
xa50bHY4hA1gCfKaDYXmfot/jGvCnD74e+NYAh2hg5JrjUUU1PJWZNf/S8LTx1Tl0AKNjegumnGS
ziLesMYi0MK9UItfYBYh6MYuJZQGaXa0VERKjFJjhV+kV97bXhAHUXuEGjyjU3XUiYjfGLDPIuxG
zqWm//UqMOIAbatgALepp8VXhQmG/BdueJ+4gb5SKe3IutiyE9kul8otOP8mU3HEoUQVn9J7EnCP
Y6qct5fzlg93yWwZPym7xMpUxtKR763GGkIxMZCBGqw05JI4QiMUZb3lwyAi9hU/4W7RvGK3qTER
LtvIiCR5STvfyUA8UVPA6wSd3oOCKU9rSP15MrM42N8ZsNWSwcMDgZl0dz0T4xZ8ZTzrvilKaBBJ
D0sIraxWh81uhM2XZiIvI6g4Gb/2bt9YYeLQSWqAqnPGJbUL4scKXl8iNwhl6a7Su9M/5pDmMIzm
Prx9yRwlSY04XTKdh8/bHYi4pIXaKHMB94TTSzJ8NFjezFSYgBQWuITCzGtqbYb7SxrdpDyOo/9+
Ws6Zk6RZX+HuGpLakcjSBaDlj+hWrdaCo91t2ljr1ajweV5GCH6B077Hgnj2SWB6Yw6ROQWuqvOw
ygRPb9qScz6lAyUuAUIRSgnVaccGb/DnDmD5ziKsGZ44T0nPSTo8tMk6xE+HMbTcJpB8RLMruii7
j1FOgyQAxv/bYY+LDJy2yXIq5tOy5jBH3NxqKR1SsnlhjZwHQqw8jdEr4sHBLhqr6rRxOo1eORzp
0ROxFc9C1pUEUJWKxr00S3F5oH/S6rxMjHsrSI8t5yVHNdbMeNjuVP84MYTdqWaOQEUr8fLfDcC/
RmgONin6LdKnyJ/lRKhWl8v16q1DHdiGQL+ZNEx2/S7COCozj53ltDPQLJrtzDJcPmXL+UnQ7TBn
fEaRjwVFZnKo13PCeYVdPY55/R262mHizhZeqUSeRUhUjV/sfgzVrkNOseWG2ADcWhIm4Lh3Wby5
8r9yCcnsk2DHHKQkMJs4ZKmWCxkEwp8uIpStvVzIOyjWgmL9TGkS99asrlo+kCfdT976CdM+u9qO
Pbr/aNaleGzdko0GqoOY8tOkmedAOumugs0RkT++DvMj6hP0U6sgmX+jYt98TLUIl7iwIVnmMf7v
SMFfs5QS/GKqLORDMKV2okKG/uQa21YZgJrQ0L8kclC1n9SgQESsbPckMmC4Ur4fH50UCIkkgVo0
bqqH5/bETOGVWU6gGb0T4bcL81ipVrARs9lGBSSn8SnBMDGYOBgHummI3+QULycn6dPbdG6zAYTG
biITlOeI6Gffn6WGHUdXXPZJon4BK64l1xu8Z+BQDYz4RsChhsT2Qt3HDCMo/heKvvdIshAZ9TD6
4F76bQf2O/fH4rRVqzphESY6sq5ISlwsL49qASnKpW4PHeIXfsezFAgzw9VXZIm/LDWb4t9japcx
3pECRIgjIK0Dy0G/BWWz+MGI3p61KaNp2Lvj+0++IIVuBxo1JneZk1zHg217suu8nUFqVyuNH7Hd
bhlzfALLMkgXF+NYP0nQkvXla9wXjFlxv9hzw2FvhadsK77FK5j6up+82/hRBvS+O4wQQMEFkb+m
kNVQ25IxORKwm9jMXuoqCnEWZqn1MeRDyua/UcUgdvEfX1vNN1tpzeH0niv1oNz2+dzT7ONC1ViG
JAYOTbIuVB+1ZSqh6Gy4cpvlqau4zeNts8T7xO8S5mR/9Wj6L7fdgxSGjDNuRHcPoBfTGsBH1xjG
yjZ1y5iWw7toiLBiSZw/GHH/VnzN0gDzeHXoQfC9DY6C/5JnfxC9KV3oyOkUdXu6LW8urTwWccAv
O+SlKrdJ3LU/roXkzKD4fQ/0BAMfl0Y/+i1jIdDy3CHSYx8TBaDBA2/1QCUKqCzVw/IaxvaY/aNA
23hF88oiqMXQ5GLn0PreUDLzezsgJpi7YCVg2xkcgYGxDD4wB7xjp8kLbYIcegncfFHM1YlYfRGh
YdjGAzyKYWXiBjI+uM6deZZe9vAyjVO7hOkEEqzywInTpVvXCdgfz+O3IZnKkhg0rDfJ9fkEVrQi
mjR1fUQxzsDr++hANCEgk9cH6J7ehdXAacY0S15tlK+wWRxFEFqxMBS6hk803oEALklytWzGpcpP
dtoRezf5ZGHlggTIjo2G4XA4u+IqKdw5dtu5lOrlCg3qJCEftpaNDl1Ic52xk8ZVEFKKpySO4Ckz
ASWetK6rkl0pz0GxT0nqQkkRhKihc4zbHTm/s1fmF4BG0uA6QuEKlUjHnXR6DhHf9+A1GO6U+nKn
3UJNZKhbCISEAdwG/bvlPM0lRvEUYEVH3kyzn/O/yy7ck1wzb43Y6XJ+2Pt7SwHYOczP/8vI5bvV
zVcRpd2WkIPDfEF/iBLfCJz/SC3LzA7NrojY61Txv3+2iohOb0wu9+Tw94vfCplJYUz3kHVqba0t
IuhS+FE/SWAhVU+Ideh2TTItSs5f2QxS+fZ588RhyFZthbthyHkQfiAfpzJ4hz7i8heAN6BwWLt5
srRHhLP/d/OcN1esm7ML1uJHndbdPxDrYe6nXGql+9DpA0O7W3yNPWdjZvmBjhgiMr/JAZiZ4WO1
TFbZhJA/VR5qVlpkX+ocDRlyZi7o/BgjR9KPKL9DBspmLAthH71im/DsPQ8d7ox3I1QL+SqLIVqz
ggzhPYfiM0le3t2yRThtemBgxme4JweU6FG186UbiOSIIMOytOtDyqtsa8SppW1xQ1WAXgmLGEag
W8D8Ze13j+Fh5QiSqO9OPlrxZGbOQRvKziWh5NZKz6W++pHTHhWnTovYowiKgXi6wvZ7y0huFmJP
JVlXewwFJrPs8l7nSLgNupaXnNJMpAaUHc1qxfAuGkQyXbKHH+jrDNb8rMuPTXbvm49s3Nk2+X5B
r9GbY8BBLKORTTBFR+PbMhl0dDCnYrzzv1J8fEZjWzdhpD8NRwhdpcMEMOyD2a86lghIp1lol3HI
TKEXFUHmN/HXhj2+CduZbRAFaldqd+XKGBjL0gK29IATzrQl1MipCeo4dTA+mZ1+qwZsUvh7vQ7+
BSSVYpNUO2P27vNUBAM1OAvGCu0je1GOQp0Ez6Yg0Qn3mWcMQ/SuLFs65+OsqpgM+ufq/PbQEdnv
jG7ZpijYWunXS7CY2RMOpbaap8E3du/8t6cvMeknyTY7pZGc1hihRLWd9L78A+IbNPpbtGr5leby
mQTD7cVJ9Xl4j1sbbBDoXGEu/NQo0UP6x9XfMiSQjxOmVmrQ9FG/5FLkPG7C8s0skMMPuzWBphpO
wPERTDs5D0x0LKVwyQa6x7Y2Z1ZQtQcRfrAjYj5KboYIRwxYEivMFm219/tUre2RetslAEFltEhg
DLBzdyibBD0ypQQ5wkVBZm6NvtuZkkVpNvDsv8ZWuMRNLnhY4nuzd9g6LkXTtCSLYD5PNIs3/vG4
+zaJhk5D/Bq4HRsUiPY8uxbzgTz9vRPEGHuxfj+kebb9oQvAifkhCCvBeqA/xGrs5xFwVljxBoe2
DA2hR0kfMZGP5mWST2qzGOIC+hsfP4gd9CTXILUlfTFn0q4dV1Skp1DdrsCTCCrhLH3bJxeLg9dN
VLw8Pc7APhDfHQk6CDYzlhGytJ0dC7bqu5o+nV/JVUpoPxiNjOwfUg3HHFCwgX7jK4jLYO57puRk
UOsJgRBlR1XYXzRFrtuiFjpOWSW40HqgT2XXQw1/vBpMnoSgmQGc7XL7cyHTCpLm1W50avs8SnFn
EKl+66fXAorCnrui3L6UhpmGDAB2LUhPFUNNmxi05w/Lbp6B/l+P8zUx/hT9hzRH1aONU5Tu8YTV
hQzeMhK0CWv9U1qOiENegrwrqoBBUAFQhKAe8abJT9GcTkDIIyO9jDUHnXNOF1CcgffpckLUa+Go
ZvZCsE01OWbnSquehW77l3zFEts9qZZUH5wbCmW4NgqUI24QRbsePn/6pD/uDdkYOU/s5xGWjwe5
oRuBI9JJ92WwWTZGDPwlTsyjsnE9YH7OzsDrHKzj1IBFPgnOXi/RIIMugHikhAXAa8QA8ijbceim
A2avs+NousHqArWyA4amSJCgQpJ7GRo/fLS6NRg5ZsF6mSYM0bSSZTrK7mrZHdiT5O5e6A+ulK5r
Qhpc8Sm5DUSM2OF3BiBXE3+Wx399sUWfGBTiAh3urAKpR+CO82dNPiLOehEiIgOZSmE+DxblmGdc
tHtPVs60ZDmLhzhUrZPoYinJpx+QVekU9Qzj5gp2Xo1e7iKkBFo8NEt2qeOnvi3CzQsx9ObsWPWR
E66F9rzT0MhAbIclRQTK3/gbMgR19pFyi5oO7EzfKCHwTcPCXSF1pyMmChIW6EFHddS7q6vwx1xE
2cGO+vE2RS27cNUc24X2rjp+hVWC7Q9MmlHvp2+67JJwFtlQ5xk98Xv9SnNDulOppdGUqFGruU6y
LdNx6lPwzUO9aR2H8kORg0k2UYbQh8EbRX/z3mOLKKrenZ5uZsp1Xa44U1urI8oEoJ82Qi7U9Bak
cDtexsRuWnVal6ksqleaF2hIXHXHgqM8wJYIqvY7ERoI5fQlHsbl9ol02MjA8RsuRjqSS2A5G5Xx
UaBye9/lCpdocWtTr2N69EmTki0gmKKk9x4nvUvXRG83yZ8qGU3KwWR4P3N/fmmvGwqrQBiSZ73k
8kSOfbUa4JcHfAk84IyPL3oigWuOGnJnVaZoDMbTDxawNXkjc7i+ECqR6auuLmhWTFHEmZe9mCji
Edl/mKRNbktoazJ1haDLvspG6+wZM7JcBAH3/xjuu0vI6sNZ4nPR0kvn0EEzGpEcGy08oWcSc9n7
JVf25ebICEc3Uptt5ckolT4LgmfVGgMxB2ZVq5GGURLOSxOt6alBNrbo3v2H1IPEIIsTzFH/PQyY
P5H6pvXjPUrZbuUU/9gCbaMfdZK0pVrv1JGDF5Ts7lOovMsfA4diRtVaOicjlQhc8UsO7zdops36
UMzvCY3iTFbhaj1uDB061lIGP99cmEVdRBzE6I1LpiPZARKf+4Ky3oz3yTKCCOOcUvsPRfoZnD35
3mJY4OVQ0PiAvNa7/z6wuPsw5/3uerd81E/TLi/MZpS1G6WXCcS4KIZqUscJATf3/RawBMrCJcew
GAYZmc2N1fhcNnVMooVuY9CdO3Bvxf9jMmcgSZO6ZB5H5SN8xCd1BxYz86d4AFqN3nziiLh+w1GU
vnQO9BGpY1Vofv5KOj1/OWd8YcvvAMkIswFpecqJ/tbrLs42hYv0eL6M8ZDbXnLEzyvqMrefkChx
vmzjByLOLdxjAyP6a1ut8MHDXutYHoTfgQ9e2Ab7/9FXk/a6XV6YIzK4l91LkgpPauGYBf0OCH/t
E2y1/hlYB7ORSbH19KcEoUJzKBrRXdSylUvENowJLxVg4vWhhxC0L5tZhu/FQRUP/7i/vv175Km6
zxkWPnUy73Ari7FIHwcwpha/Sqm+O12ZeGx2BY5ytya8N/0s/qNOH2DLNZPJ9JztQziskxZkPr6p
cIv27vYHsrF2SOxD34cVFFZBg/+in/l4KXrS7g+0/pdfrXc93x7wnPsIjvoAX8DbiixtCIq4I268
4Wy/aUvyd91jFobFOyBLQojxD9oDG+fKoW4auQLvjRWkeJ1BLZnEskDWrvQOa5WBbdgiF+2Ts4V3
1u4o0R+m7I2u1keDRu1nnC9H3IhoFmUp35LsGoTj9Hi9cDcDFjk243OBcbg/YSaGpEAIkgWYuBKw
OsZtM1J3FDlMpyJJL4DTds3Qe5uhjF1zlpazDFsFF0Rojp0kUm3zgdEzPRk0eSfD7BGv71EB3V57
xLW3bSSeOjmlxEaSRPU8V0tUdiGUJpQNjjanCB7d1yFlFVcbSNvBdavQ9lwXKgz3HwEfr9Ptbn+b
ytd8CEAnYkDjkmxT3EI4G4mijIWGOCA82oBw0lmZ66dxa2MjL80UxmyjoZjkl3e1Wyjq2YHBE0ZJ
R0d+73oyncso4cK2xv6k6AX9JQPNiHZtAB50uGQ6T/eOLFFHXcDvsgoTiY4qXbpml9HmRdfFaQle
B7mbpzbJjkk5YaCDs9SGtNIYbEEzXfuGz2tjJv71Du+/FJGyT2MFUmZ61HPHCQd1B8KGAEsO+xDv
wlhYS2/xoDYead8aiobcjbCDHnvnBJflQ3DUkFJpaxDT25oSzCYlBCjF7q/mk/zBtw3d2fYDPzfG
S3K7M2Fesu71Ne2HxS9TEsppb9R5qev5I/ibTgkbfo54vMU24030D8Rf2xlA4A5iOAWMKnunR2Ce
7miHjkyxM9L79AM6Ap9mDW4JCGWAzXb49hX+pJGHMktYrUV6Tqg4vDOoxin9KZqE2E+64+Int/bo
0/u/n4147pNM9GAYhbjFOtsn64vqdLTaTNAtJQgLFzjm7AeLDOQMpkU950VXVdAep/leKyF3xELP
1jnXtNgpY0rplo5chQtrXbS9WmTbsNNFhsbYw2wH+ZliuDE6srsH5mh1yzMo9jGS6VR5Pa4m3NoD
ANTJj4O7LLtVJgo7alFekrQ+oQwPwXdeyUbWg8E78JYyjDkl0DBagH8MELy9FkGF+K0m+2/DDvbH
fa0C3dFwYiw5yQao4SJK7R0+c3f95q2ny6c61ETz+dwBRbaKtZWDYMcYFmf+/mTyuEJFi03UXqv2
wi/k4E3AJpPBibz4sQVic0a5zkS4KRsHP7YgzojXrsbf/j07kC1GqJ2GhXQwT1DmmfcXLGq1G/qo
LS0iYYSuGZyMkY+xgnrkCdPVIrq5IEtijufnZDWvejUmGRJBowIVqmO/6fnXXaN8Zq0UA36xZMTq
NwD/hfRcXRMnQj8ZCSa3EVX3kAYdUmG97CO3QiriSvZyeW9eQuCnpaFEYWncIHB3A1UEyzB2eUhv
F4hdRZapL8LP4koO847pdWnEdR2kZ9qU0Ka+Nt6/VgMOlj71bCRu9rkYkptwElzZqsQ/bENCxEDx
YBNciPtYd2fARpoOYYfCLGrwuME0Egf27KgPUc/pbuGzsoCaxfiIArVmWXev5rHdobJNkkXhbKGL
xUQf0OM4q5L40Z7K9c6eGPHTD/1gqwImmhtsZVx8trrGMvabyTxo04xnLjUIkm8SMn31WfsG5ovP
bJe5rijcqRpakmW2iWRRJTo6jJF+XWqFL+EVJztLpY3XtdiqlGmEo0Bqs42u/gC5UOX8MV1Pb/Fh
jvDJexYGELJGPu9evfVwGMzypYot0mmLlbfF1CcPIcdqP7PUl9tSejplHBWRhYZB0Ymn5qHCIX44
WX2lu5wXfUWt2TnVUQEdSF9BdIlyo88CjKeC1axaTWGp3FA/M94i+MwluH1QScCdPTjWWHK1mLL5
Q8KbuQJlsxUI5eSM428K+D6ZQ4uzjb+V9UpnR+BuKitT/QjvxZ3yUfoF6+KbXs4Zk2/rK76h/INK
fAaC3MylnkIuq0ea5BKTHck4NDLf/icindpxiSl8SzUxVN8zdqMfNDzGJf4a49s7WSCmyylZRG4P
QLYJdlJDTaR+pW+EbeFsZLEHfNgZsnqbBWgNDjnXBqvrbqnycvQpLoDOBekoHuU8zHUUr8Q14gY0
BEjRRjRHO6fE7SIZbjD2zh2xY+43HhTa095CnE3YqtyK5oovHA+3dJtMb7JVlScgsK/tVB6tScEp
COBm8TWoNTIrqjd+HKW7peEYJCpvFJShzNY/yV/0VqoxCwSScPGO3SjYQkj5ciKdeLtP3LXfY2E6
F3je/OZStLQhkXATwoR3zKZIG8pU3TL9bLCW3578pZmB86/RaiFpb08QG8BevfRoCPlvBGpKINK/
44H+cw5HgkFa8JzS2LQ026UaQNDcu3tQWbeTvI08oODa3ZzXlt14Uz+oLMTumDxNE/Mw+I48piOb
D6k/8/Ysa7iTWSXHlAwvgukGTOit/rnTlPR/ErrClEscj7nrfbnaUk3JH4Dj9SAyvgrySLqo4oVf
krrJz7wvYU+bjGq2ilM43M1pUC3QbTz1kPq9RgBoM4G0etJPAzFcj9+j7OoZFJbDo3PUeY1HfHN4
X88lr4wYSbjHIaRC0bmDZoukMPkdYecSw9oufxuFLpOI6uZ4IZVmnUlNv6YtBoPqtIW8E6zhl0mW
ikfU0iKHQHWlF/bUNpZFX5ZXsnROarouIJQ9VvaBpOyue+d61Yvzfb9mP1T5oOLwlEMfu/yTVw7T
iByJQxD4+lcacyuajxK3O245gzFn01C0mBx8GMvf0IP1a4f3LSsnAo9Ew5816QIS1BLUfQbWJAMA
GYOtIrhASca25CBH2j3Up5kZORygq5fIiUsKcm/AI1pR6xakNYZcFUz260+IAsXLRL+3ppNouF7/
tI5ut4CDmQ+icl5kVOK1K7YYlkt307rY7W93IqcTJfuGMBaFR3SFtcA6lPXvkWk14aLPF1fe8z6p
TZSMWv22+33M3Fdl4TLXIE3UFdm7Pq7eG9UGnZLmYX2h1dCsE2ilL6/tXjDTjTWO+ue83cYPoxBj
pYIpti9Q24h1itnAxusDVKadKzAiFQdyvmSPMnp8dww3rKirkRhQEPrLpc1H5ifq03Cgf3rCpd92
g+7m4BWfWKSrmyapO2jRMy2r4LNnehxCc1EImVTfryH9SnnC4RjPt4l0YfzyxKCpPml6i9iVonlu
3JgkabndBmLp+kZ1gjYvmevzz8ryq/PLcJnejKPTHVjc5ZDHacD5BSckAOVnQAO/kscQ9mO6+0Ld
rMTPOmN+o3yms6D6qPTqbvO2I2s+xgjy27OeMIGucnHx+/OU2esoNXTpUYOIzgnYhsh42PIif1SK
Kn83BhwK1mcVdTCET6Y6pt+KHH84I9dmC4w5Zhhgs3byj1L9HbiZ/HPBYlnXxuPPuyBoQq/taXoy
h6M0jDBy8mBB0bY9afnj9zVtuugjoB//ewuhoipxpPb0sd8Its7/jigPQfaFnpmyw2mLFsya9jQG
kv11aJQXgb1aFhKtWukDHyJS6fgK/vSYumlXWsTcrozlK1wuzXUGgQWAb3fCU2gUGh2hs7E5VjwS
At3xb1mboDHcQ4Uj7WwPcvB2R/etFkiNSzOEbeocA+0ZAL4/kyTBUCxvE1gmWbbbWO1pxOIMNjaX
VftaAy/Zd9t9TQcvjom69545C4BfhaTwKfEUfQ4ITp5pxvF4PhbbIRY++ccy51T/24lY2MfaDSVP
f+pQkZJs2ZauhHqRbvj5uv7nYmNlpdMayjdH37jRksATw4b6M29QWkKhG2iI59fmyfLp4BQpArgb
kiGaXDUEsHypBI2K1GEWPwjZKyo5+lPR1JmpZnWjORmlkAPM4G+ObxPtDqz/lxhHqKe6sPCK7Dgc
LRUJttdxqeRxOJCTEJzXGZqBrouE6ueg9q0didpiSqmwDKUB7dlH1JEIMZwwm4Do+g5tMRkUkzG1
sX1MQynuXYlKLWWxL72YCnLdFAJYkE/1GLIiJ5sTYRoC6qrq2RHJMJiIMnwMEUvYenoFhfzeYTxF
f4BD8rA3YC51NdpCCaX7aHtCnBj06LMoe2ky5LCIKR3jo0wh/QKtn8uUGC+WtDYxjqI8rlOGBezL
Nxj5OlQsISUQ6AxHLPuiFvObR3YUX8cVxezfjmldjj5OvpLzhiM6Q/vDJFqWwAednykuDVS9WH/h
0xlt6UgABCPVxpXV+akPF1CLd7lcdaxZYi5LLgHtijaCZ44zpPKXphE7d5YPBmLAfNdNav3o2WhA
Vmtip20dvJ5vIhxyrp7YZM0WcBrIZ8/cyHKPq2dTf7hqn4CshIQYs5x1AE6Crzj+3HMAPd1LN1el
fTFJI+sARp6vbreZaDjjN5q4I7+3lZ8S8dYPv25OTVe+9B81cq2UoeZ3WznPrtWhDomjJNZjLypr
YrtwGhvJT0rpvVhwP7HmFdEUZiiIDvsWTk+QLBYOBAV4gGgYAedM/PuIQOhgI3UXgposyf3vYPqm
qTkKzvfymnFC5z/hv7C8klQrebs8Tg0pIO1/A8XLQ0oR57HzK3qKams6fVEJnLTo2vwxHqIhoIvF
u29XSvYwUlKIYJ8uGfdl5TtTARCEFrSgatdzoCEk5LKCUU36etnye7SzRQHHLuZHSoKWBuW9zyOt
HkAYWDy26qbo2MnhBDN/lURw+qiapkUIyAu1+7B+a99eb5DjkdYTeCQF5U1ymW8dK1hOdTc/o7xQ
rZf2OR1iiYKhheEQfM9RqM6L0shsNiWPFANZdeISYRs7ewtzuzo9NjF4SbeQIt1d7KJA5126jzCA
rHvWq8B6IwUxavG1Ur+Xo+jmjxXQdiGyTlX/WodGRDDV0LyrKv+6ROkSUVuEivdEGQvi5oIL7btY
dpNGBknBA9omZuyrWvgNXHTtqb6rFjslphhrwARmWrOyE45B+vXfD12oj3AtuSrW6niDMYmLNDyu
srv6ceTbInSy2mq7AX6zCzTav+rUzWGoWBYM3FMxha8VbsY4DszySJWIn6OfSlG1ZJYb0/3Y4hKC
4t/dC6aE/RlVQLK54Qo3froLTG4gaNJW/iQ9OKPubunYVr2xz5AtS6u5AZiR94RPjWOlyh7KG6Vi
UcIxhRu/ceyswb0TjwitNY57mJi2J0VgzoQy8oOGP4LzHRgtiBp8MS2MvWLVJzqGbGgyYn2Sfc6N
hgzTNwSC4Ko7n9cioTab2VYObhed2EQbRpc2RI2uRmBmrRGOFZIG29e7xjrxDozzHCheYvwlZ9/u
wqtrFKQoZs2tnp4rTydHBWSwlUdYEO168zjEnz0p/35wYfLBorJIO1ZMjQxDhwN6h+nM/Xr0vRBH
/BgIlE7AthUXMY0kO2+bmwH0iVf4RS08zl8uM0pAa6L8DD3AwpNHeZuyDLMu5KCtxKcBkcQvfd9Q
dBmM0YD+rxtkPgwTZVnaZBSLk/hHJ/1QP3JnnoCOlMfDuiUNUe07htYRP0Y/kkRFt41YWkJY45fI
VI0J9T9CdU783dJxjNCZJ47gO1tMuA1Hnu/tRX3E2a3x27AOfb+JFhevWkkbpVpmoWriqEKe/Oxj
XXuLdmI0qoJWil9Tme18hgnzBRr2iVAxK7tArI5iejZLqd4GUzKgD87n7/XntoODKWz4z75/6vOr
CLAGJdJdw5wORDuI+3SIb8XXI8FsuY7OzvRKwzMsRJMH276P7+hHmPDf0mqUHlVH1NgPbsbcTFos
L3vny/mIM+XSV7l959Byn4+aDfpk+nllFXF7mik9kEUExFIeK6TMApekYalz7z5BhCrdDjVWKxgY
u/uZ/e3KYoBjryxJLeZh1N81/nwg5LlqC1hCM5HQ88kdHIAfZLdNAdzyxEcgMH1CQvsn20RkJqFz
6ohY3xQ+N0kQyjMqNs+7mkZgil/wLEBGMysuPKi8S9z8IEj86KdmOQQgupUQuYaynnkRRoLm0xuK
W0a4UYjpksbZzylkrbczurx8LbBkAzKYbe++RGiW63+FmNveaL9fmGCbcO+JaQbzlrt3jjDB0xHX
H00+CNzq6S6rMHpenpUpRKv6CnuuYYfWIA54htciqNFt70TVDvu6jqUTdAYaKe9yx9JTOXxXkLMn
DWmCvclGtcm66JXj7XKV3qpoFG8Bgpg6s3JUqrKEBy9yI0gZQ51EaPr1YHWnPewkAni8k1QeXoo2
iv6ZUfvYBENQtEfDJXgDD248+L3g3o7zW5Fy9sp6sfO+TU5A9OCplZCL9IiQ9oEmsr+fHVPLFyTp
f6ChwScOD30HE3m7iup+RXB5egks2othUJyKewHenNhBvLjkBnvry23dQPlskvxO3CoyAaAXNDsQ
cCt6fJ5giX+jkqHpeHSDm/K1cplO9XHm1s+VzoV6R6X6E6qGIplZKkSLgS90J4W6mOQiQJenJtqT
CwYQbyzi/1PuOleRgKWYqXcFQNMqejMqgFZuQ8Y5OhvWExsmIth5VUlr73iFPpDzwH7+FG99vbO4
ogiKltkNmLTQ69vTLppp5cG3Cqh8Hb1uX9SJojxZlJQ9UOyr4bjBwtkmUSSM2yNqtvhlIY8UKcw6
5UAU9H+5Cpv3dLatRsgkgGWqphzYXIAo52margUF+P7fwm0xrbHqCGiLxY6Yp9MraLXUTdgoSewi
zh4oKtp3bsbZa7KtfJIyabUUl9zgq83rwN6kP65p0NSJjNWe39GCMzk+7RH3yxGq+fLR1VleipwL
FgeGkC0DgEoxt2JSastJWmNrzGZMhpnSfORDw/Cnaoh+r8Puqop80ZQQP16BvHQVnpPBoqtM5MBV
sHhtZ33oQwcJn5UJ+M2OgrLKC/G/rg55VKxgBYfH7YIkne4sD5SleLaN6SJgCAx+Iy05YLV/YqhQ
56lPv2QfIMPQxcLgEOO9evlHPDeo3YuDK8O25eAZniaC4BaVDFrzNmRQvwkwvniq+azF4cALJM/x
rkRIeyqzQ44eZHx15th6iVfSWnuj99vKnFG949IIeJQ0uo9A9V0MxgrvsPXIW5NSriDjd7RrTaPL
/yKUsBq9/fuyC6adxXcDV/z/1npv7jG/8SRdhHCQJEzC0Rfbu+J7CGIWaSqTyBNMCjwQAgx+EUZK
ktuGFbeioCr/4iGxOjrgoC41BIoiHaMuvy/Ja57jK32snPmj57HfUKgmewuVN3izA8ynflOmqhaF
g7PN+1I7Xnl69dV8vtaVvb4xsSZvrlHhF6XExsiMdM5W21BhMr/tQ2r1HNdIaN0LdRym7TDJN1wk
E0mVuKo42Pp539UDjKA093m5yWD702A7rWKAvG4x7I+UMKONBC/YhAE5uQuzy9MMSRt4/+MC0ltM
+HXrBP6bgwXtlpsxtY/fM0OfWfcm7ldVW+AO2FA4KlnIQUPomKXOUlOhslwC463Qsj7uBDb/8/zJ
XJPHQPVYUXiQBysPtkeX91+kavnSNGWOWplj6RpwQMC/QCV5FeVMykl1UY1dbCik76ReMHdX56TD
CtRWe6mEnIdWmaHHxpgLmLm6eB4MzdzLqzHbXZ2FtDKnqnLw1Tagd1AL9tJCjDSomkwvIDWThbPr
+7xrESAlpP0pQp8F2U5NxQcud0Cl1wWCs1+kPGugGtRYrvdWtvMS+gU1lk2bKN7UjmD9IN2MEGji
FHK7YI2DxOrw6ELJBJJHr6pb7YLjaYUzR6R/8Jq83mi8hJuN1Xl/P+fJf3KQBehgVqS0aSsqQCnF
f9/0GV6iZxCP5/fPjiMa/JYmxBJv2owBrswltjbpCfWhcOgQcxCOplcr9DwSebW57dU7slINbILh
NcB3aTPyGFaDGV2C73fBmp1jeJu4BDo0M1aUcr6Y49PmK+TWDCxfG1bNXbzUgaBA0nmVZseBYEtP
lvjDGT7DT/BOnT2EudvVPKtgLeS/sGBOjzG8zPA60Ts1dwX6uXY9FSBQ63+qEpZDDAwXty9r1g98
jw0MUhCPT81IPcdcKccCEdRq4PCsE/eBBumNI2w8Smus38LY4S7AxQEpnB6VZclqTLtfpI+ifUn4
z6a/WuQwQ2CDV37yZtkZfA1k9Ag2aL3yjgjSdR29zF7lJu7TN9Mluf9OMSnlcjL/l+QZlvhesPLW
kzP+kbNPWPbMYWVhpnmsSmtWwAGGnaUljfNC+0pA02+vP1lfWlLV+77fN6qbS++iU91ilxvao13x
4FXyEu6Ftj9/shXhPxmpJSLliY8MvLtU4E9fzDYNVL4QZPdPLRPxE+r7gk2NJG5nMK8dWVTodfVD
6ga0O66SFBIy2l+WQfe1HyQVEXyu/QCgf+xlTaSolUqn8lEaavrOtjp04D7EvMBxUWDFYebApQrK
7kAtc2nZuz+rPcM5/JX6ppcWb3+ylAYxAuaTTEAp0p+b/wsb+iESJBuIVsKi7f/Y0IinYfULSgG6
r3+nAY+UEgc5r/vBeQCrqvRVWh14zRYqFWkwMI1zJOldgCo8saYL2Pl8j/oM1eTI9hd4fW7R0s/Z
HD6l9R+Th9Fi+xRWMWQbFhdmfRaQVTf/iExaxtkTTRcRZMExuPZDUbHg9JpFaNlDGN3L8YmIcZfB
5TI4n4VQInPBfCaIJrkJ6cG6vZnQTy4AAvompa7mP3LhryeTvJ+kB+0IkiTgzO9WBD0k67rreMuo
2XuDipFAy+TC3c0lAFBOj2bEdIQkRT8GqmLMT9Sdry/8SYvPvZ5/1q1TXfAFyQUxTMqyqokbj0Qm
2ZEX4sEd722qmp77x4SWz4x84gsSRNEOoaI2x+oFR7i3KaV9+6NIMb3kSC0ftbYXq/03c0ZKDUmo
AwQO47+kusolLHKdFGXuP/RjYHxaHjQ0xiMX+pMV8sr6z0bPpg4Wmf6ViBD+hqlFdlnNP1rqPJz2
wzL/R1SHr1bw9ExFJ7pvVPvCVqXtHCVd5iuw2dZ5/pmefjb4BkO2CIytCYtohBt2+LQWHnaHMW6f
ddCRlteiOqvdV9AAboqDeq7WQRbb9MyLTsuKixEqrnuQlMnDIyMGOeRh80e0qyR9z38JueS1u77/
aur5TcA7+AuUzIsbbGtis6PO7tBwSk+BLbUx7dMC2Nok4HjIMjiUxXvkTReVK+mKPcS+dYz3mWGb
KS1kNbF75rHS4zUr8NKRssKaoi82swl6Gtk5RA+ZZcgJ/kf3oLr6EV4rf+0rkfWUM7/ATFlA04nQ
+/TPzMa77wQs+MZ7AN0tQSVuQnLmLAwyXWRKjJbISy9uKNh6ZGC8CjNw2CrDgXA8t70Cm5lIJq42
SJ4CLPSMh9ZJrDl2AUEnOC7rXi8l/Y96DtI3FqkPNTPYd+fYrT23sC1aEKB95z8FgjzCZdyhfnTx
+6eGv+T5HgWDXFTUr9UDrsUn9BwQS4hjTwJAL4ED3DD7qFRKBA0A7+6qbD3xmb338h+7UK5Jl4YF
dkmadayoB+i2c0pr2EGS7YNzsas4mTtN9jkthNnSceiuqi4qgQGSQoANX2Cr2pV6tRazMfRCZexX
/pWGOLwv9ARs6dkhknw01jHQZnkOKLDZx5QKI3HeIq9owW7DT1Yk7xGF+e/XYPRaRmUCno6enoM8
/BhSqVSJE1c1bGUt1U0I2XAgyn3vnQA0ew9k3DtFkNBVZuyyL2Q77qMwYBdXV2YfSJSYeyJzBufi
2FP7gA4g96eRgfidlMu5bVSnLYBHfxllZJXpq0qKt6lQkC6YMh/9GOSnDoxxh++ud82juwAJEgxy
1xpZlhPq51d22VP6Cw+O87wIO43E3KLX2LkyzhswE68NwF5AyHwDK9B7ZNB3AWr18Epa0x4b08WP
vZgrCMfTRaXBV+TE3PqOy6/e00i+gWm2OYMQ/f2j/5lxipvKma8uNGoS1jRb25gLrByTFRvjOaux
tQO0tzWMq2FJ+OIg8s4jDLQuecmL/Wj/82qe1gw+2TAYR/Rfh6x4SqxE+3e4Iah5nGYXgCINBwSb
MCBihK1QYdvZ6LgpYeto0aHeby6gmDDysMnW55Sy2mq3flLnr8rNqBaHf+9zYXlrMCgcK43Cxm30
SrsDCpzj6PbsgXGNNYLuqpH8FoDNfHW3Tu0KUn4wYbrOh01LSJpYMLdT/Ou+RYTnNxiXqVKHuokG
gwTiov8cUvF7sZnhmXEpex7rujnQluiLYI68FLnoW6RJqh/qiLOCS+sq4aLwC3wnrPVscialvRvH
yhNbzULgBbwzQCbYGrHO9XsN9/XfmLYoLSzJuIMo2LGWAjZiJmTGUcTpGVPSywIyKT4N3YLLfWGv
rz8LYY0TAHt+7AubZLPOcTbYT5hbkg6CLvPASI5/N7q+yVevmKdRpv596j3SU6oxcEl5Sh4a68ep
7rMWJhjYyP70wD58zXmmhbkQ7IXMJWar1Ga93IfOuQxHQeAbtjtUp5P71Z8ClpDLbxbkLlCpllMz
CEeAVtQFVbpE+NpyZhFFFjCKx2CrkSN1KKNL0g5Z3PGXNhOmKR2bFKr4YCMNRUV3HWx3iMkEPUbW
QVmOwJs7rPOr2QmQhLbk6fSTw2/GJVvPQXBO6T3lTioQX6Y2BL1eFmLu8d/0PLGgTExSU2KFhDxM
B7Ee2aigE3iGUEtxC9T/LJaoZnA612cHojesau/ovUz41MUCSkWQkkrwIfB+K4dQhlgxDeD55Dnu
TJ8T0/TCJYRsfCyLH5m3e7+kK7YNPHq4tc9cifUDz5MmUoT5JkY5dZtGnLexiKdo6sWSAyaAx9iw
ihyOsdj8AkT5hA6oPjBezkRuzyr/4btOZPrWb0DUD2Bcwg2K2c90UZb4RIY4WjZmUSvMT9afQZld
kZ207PqBKIlB22wq38KBnxSdi+I8G8C7lEnVlAwSQBeiNWd3M+pudQK5Y52eo/IOBvXISRYMAK/D
lqIrU3t4aW5RAqKY04v0/vFmFYMox++pvch2dbg8i+1CB7OPWhRIAKfbcPZTfMRaJPE0GZnh0wdW
I/6NflVGcSGui0bMYsm/ieASm1bxOGRq2XwYHpbw8eUBF3LKHGjP/Lj5haev13qGhbG6POp3iAQF
p6pB1XzCFEQrwZnNFFA7BFsnBheaN/mpXJT8O7bcoC/EIf+YuQTH8a5hHJgcuFB5tuPFzJGu2C2i
EK64RC2z0rP9gHdVcF6xAQxQk6+Q9r4cMBaMlMyuGaOzE5udFh1FJPjmZzGm/6f6SeOlfgaFyx4E
Sw1y/724KwX9AqPOrWaofRWZTmbU4xUhFsYiplgGmdcRDEWe8gdoOV0eztYbDN4r6r8dEtl8OTmp
9GjPr34k7PI3F58ef4XcOMYn0UKdIWMCqRpGOukP5yI8NTu8NQZhHD4AJv+T4SUvD02aGbKLOY5D
fvFzM0WlZ2F4Yn3yEFv4IgzfARTaEZBvni62ywgoNSYZocCht/M4U7dM0ECwazuZkeGv6PnpIhYw
ThPgd6mwCooNv3aWhh7Xb+swAld8v2wZ/Z0hvgzitG7MCWJGSzi3ESqZXY2v00xT7S/bsL7uyCVo
gbnjQ9k/G16KT4zzFsYvRIyjc3xIdYm+dNfYFfOTbWkWCTXfPdOAIkQBXaZhgKd+ryKOdNYb5qAq
bnpsk4uj2BhtfbAejU2jckYNOYz8183RWEP2ex22glxD9ygg2dGeTOyzfWY8F+OeC1Vlblt1g7xl
TdH/DkwSavng0fqK7OY0qFkaNmr+u3SA5DAbjwXufVGawVUW3Rsur22jOh75F5KjOhFj79sQb38d
9VqFrRfCfPipehTzTTufHPIrmY0hS33012/4yQT31BBuL+QViaJ5XIuQalYALjR3J9y/o52vzZLG
C+DG9NfJbwU3/czCLdHQ7+Xlq//GvRb41uyVS+hdxEvQ/5NTlCPOiyTWGD4D3lBjirVayLwBAIc1
b9qdQ+uE4GGfpvF0SOUb0KZv4n2dnOmszdddYh4qE9awJhvi7u5KpgM+AUOlR29YZxTYjN2wgnog
r8miMVkLzzVe5NbJLTZWlZMDt0Kcj8o8eKOgtYpCCAB9Amn9vsZ23Oq0svRucOM1bFdP1/z0cw7w
Jgr9CIc1zd1B1mIeOkNucI9AcyPukr9ey/Eks514wTOI4jZxSMHxzmDNph1JmegQJobU/05HBbOv
TJU4wENAKOnpf9WPLe1R9OhRa4DATBFIvwhgJjP8SGf0cRvXRPgfsZqHCIlh50tIWL0KJPxeOCjR
hbOFYNF7imWwBP+wFBiMJq1iqhIklZn5bdYp0OuSaGFbT0aa0ShycmC6GULGurBHRtf6zXGxJc84
3cpzFpVdlLad/1jx9seXdFYKoA0kvjV4B3gKDhtZbBvQFFw7DOJVWLNt+/vIy1mlCthq1WBrl7Ov
NCPwKFQByKVfeJD58c7Fi9dOQdvR/a2RkzKmPXhvNphIaHpwlwm3aig67xN9cAbQYds/w60ubYOM
h8GrEfsK9PTwlWLtqyuV3Id6D+CkmXq55d/sJTIbXn8fpJ+CVaZ+3m/cw1+wIDg+yPJzNs59cLDC
4juJWf4h04N84he4BwCuwTgJZ+jlPb6oohGhTniL6dx0olsMTQHS2Y4QPtt8d3ZmZMeXxYPa6DHy
wujGbaUiEAOMN4Yo3FjL8PP57wBMPBjwhP7RslJdCkiajS7TgYCVZ/l1Hak7+QL941TXDLwP9Zf/
21NTgLqTVcSgN4GPeGFPkX0WlkG6tSkKe/Nuw+927hf+EEM3sLe4V1ZK1eRiS4XN7s1g2GpynR2I
mEewOiE24hKsRFr7pD2nn75zqrSae8rBZfFb8+OFGOdUXyQ25qq0lb9iPgMTJh5q6kUccw2GujOo
Yl0ckVYSTIFgTmV+2d6nGK37aLOaXX84JCIcgTZgc9H4J4kKUZliOcUHG4Y9tFrb2busANoUe4+S
NydyVZu7Hay0jh31sPqSPwU4JqxRtAzOzSYnq7KPelLYZ6zEFvK5AwPXktTyBF7VGdtL9B10CHHG
cQCjE81m7dNTSHivDAoufcaeGfdvfeOQfrp8+U/llr2kGHYOn9Y8xZy0cbSiCXOtR5CnYGWRXpfC
ifSjiVVXbEQURojdxJMpolKCHFHwgNz0WI0uiAWvY97GhwlZhRVHKWYqc+oyi1QM4xxxowiIMLgS
EmpimAg6mxiPpnah806geBp2ENIjwBxHUiabSqtVDR0sbsVIpjZOlSAyqOdctV2KuHtiRAZOQyl4
QaYD8mMFaYwweb/LIVTXNERrsdgakHeymDE/z43WO5ZY6It2zzocprOjDPITBXABbU/lHR6xdQkZ
06nUpjEmyvwTeDIHcjmodIgRULNMt2NJ0c/HUoJN5S2+LsUjDAzt29Nyzi+I+LkRPcuUYY/bFnqU
tNIgT3W4V1azhanfZh1qkmMlzKBiLNUJTzLBfMfW4ZjOGRC9nsrflhFIqreyRWQv4USDfdfBoHYY
8JK/tGseSepI7L/qMlbKsVRsHntr1uk2lyEpM0LRO+eNbWUdKjSu9I4GREVm6FiLoyDCmWx7GLjW
0/zhYDrtJeJgAQkiuf6a4O+YPf6C2p7DqV+cOyB4zQf/l0V625RkPQXq7AwXQSOJoH8yLUgsw5OZ
saDQY8xSV1LsRKVn1uGq3njtAu13kl5uZYVN3wnBgXOUPZX4FF7RnCq05NtEj6AQBIC8rKJFao9S
2wbvYnrZM/EnjJpe2/gPM3mJ8Zu6TzbkUx6c6s+tQFN4nDZ9XE9ZZyobJXB6C9G6ny+Bab0Vsx8X
nROuLnvIJP8InskxGJuRKlKa95VFJNoUKuSqYv0YdgsetMtVoVDOAdZKsvtvBjAz7D7bVsZIl64C
uJWQhRGXgvbHw7Rf8CoJ6h3Gd0lwxoeosNVVHQ+7z9Pus+2L6DE8utLBFIU4MygDLSEeR2Nbktga
MqjCjg/+B+aSeqX1idm78xH06gHi401rjQACzrUd1catzNXPmFG5DhD5a2IEQCmZeDRaep7b3Eye
W3AwuC/JsXi1YQp0Z+qVz6CAQ5mbO2bvY6PELkydq8715GkPjjfzbNuKnl0HGI4XQ2ziWFAwQGQr
UVlxk3TXVnrRUkJEAsfDpEWE58dEglyV5q2tP+/HnS+Tq7xI6EvasoB21/Mi6BELMQKAl5Wf+rKo
LEwJcdors26RVBRy4tQGZiuyeuGEcH0v1LTJ9kyFIgRVdKa9LzSvoYA32Nodk9ropt2LWaqAAptx
zW8aIHE90B/lY1JA6vnq79iuECOdtgKUH458NkVOlox995d9368sOznYxVnYFthXFQrPkJEHqU/I
VCFlvsxFiYFqpumfXH5xJ3HRde9tgRTb8Cbeldhgy+0c/vtdHWkLaxmKIdmeFQErDpFjbvRcdzkV
4I5RKpD0XbO3B9Kt9dL5mhr5Y5KtEkeloHhU+ZxF3kD1TtX9dpT6D4sIg0M03+qaaNvNg85qNMmd
4+37PQhtX2di+L/n0n6wz6m0VJX7oiybn5sEGMPtQaohbNQWWaSQPQAYRCQ1lTdfeUWnXee5Ij8w
CD4GQE+BzWVhGN75zpcFXvbgxJnbXOa0/MmwJ5B/Qo05cS0tuHnnzELdly0xa75hFgGZXkVUu4Xo
TLE0o2vbRaJo9zRjQehuSZooWfVpTUVgN0cK+5YGMjIMB+8PvAeKTDVHtKIAlpXfRJHBHoimECaQ
OYHOqMrZDesfgDU8GyWqM+UcH9sKZF+AfO5ETsTGpXCEWLj6WHenx03copO2gGwZzFh35cxziw7p
ts6A0KDZZhxM6Ob4wWxESZs4FzOom+7bqSY3589bI+lBZBeAYcTS44luFy0JirLW3uNiS5H8XnLM
0SpsVFjKHq5wIFkTpFi3wj1irDVIaZtyhMcjMYkTsKwlMxcDd3TEz2qnT2Z/tweJ2EJtAuGgcbQF
TlNH9krAzJyNKT7lnVwpag5iLj71kn4UdC423NbAVwHknxqXI3a23su8EQMZyUIf03t0UNoR5ejk
erCY0XUlnA8oOPOVL1Su6yjFVC1za0bEC0FQD6Hk1LFz+GJXOC3jfmIbvhHy9nfmNoo27fcKIS0p
ZO8TG6Gs+V7xjOO00GWEIdyG9/ouU9o63js6DBoiTm4TDXpT25EfLS9xbERzD08ED0Z1rrwprOwq
HUlY8/BSddjy6ZmLNM7AnOWZINjsmYrTESqN5Gb1Gb/9a7FZ4n2A3dw4J1Ijm/3viF7CEmm0KgI1
5XnFvwcs1zi0xSJ1Cl+3x2HJB1sgC+cKMziITMxhmpHxfxVDOjR7KYxzM0/h61oCYuXvBIfa6K4+
eUdXcTWUQD6zcwxyP5O9GtJWy848PIOcAlMxa6umAs+BWO1eCt631vsdDpIpo3rr0q1PuTMpeCAC
LCey+kyxyAXjpmLG36geyMpfiHvRUNksumePzlz8GUapHQcMM8MkZ0VuH0OkcSNkeJ3PDluAUGHp
Dxpv4FvJUL6IDDi9JW0f5/bdaKU3HksuxtFUqNuNHJNULF4zJ2LCDP5F86sMUtO8XwhuTmU7qcF2
GGtqil9WswYKvSiQCHSpWUeXgPxX1R/Ix/lOLsfekgvxZn8uTXpw64OSs1pGFUZHiYEMXHsZRoL/
C/MOS+wEp2avlpdnNLQhmd1Fw4Zp+T2UT4LCKt9GEO8lufs5ruI+vJAVC5hJpNxxWuNR5qjQJM6h
qR+I8cLZ2OpohJJKTW2eEvnq1FxpGv7vuLQt0u6irfNy+DjsyYjUfeZwgk6JaALC4JVrlF3J1fUv
2RNqqOVW6w00FnkMbFuPbjKJriHZZ10W4/ZMhlIFxQhYSj5WWvorpuWJ+2DVbBwIDXzL1uftT2cA
3K72FIvxK2SGjlfbIUzyAX9c3lecJC9JxiGYnKOOOFXDGsVO+HYqYaTi03dTGVr9u7adSdgF2VMD
BJTFgA3/mOj6mQ3PXYCjQwUAX/FqrvxigfwRJFTEobgsq1BKakZPt9JzSTIXDI7gsi6c5Ep7FrkD
oGOwSflVuxT1moPtNsPAMTKOWB98JNOLxiQtscS0yjpXrWgLo3PbPb9ag3RqY5jT7r9eZ6kh8u5p
tT2X2iTx6X9b8AhHRyxtd1yP746uBRX+O4r3DmoGA/ysqqOIYiaQFAPyUxyZgR8EaCbjWENdFIVg
GMYnnrafZLoAaqzMtdPzLnCt9RcYp+s+A2Gej/mMZeO6yZG+WwdtAhoIu39qThDANIc0rVG1wg0J
JHYkepC9+4U0RzYhoxWzVR9e8NsTUdZO/KeniPTOfpfem0QvSQ+rW+FoLO/J9mm2zxlMnz0CHdFW
f5uW6AqWPYBQG0SBpMJjcSH2swos/10/cEUe6hcNAndfvK2FUzlJQLlE8TVxJ5RjQdL6hF/gd447
f5Xtrg0Ef9bhpwYutlbXO9kJ9N7d1TLuIp6HJswBuCER4006KUDbLMKWW0JCRbXBrZ5+7+tgqUvB
11tfeHFxv78bWCgvRuzZXJpm2U9JZO87SA1FGP99acn+9ikaDRKsCnFy0Bqq8Q1oTfPJow07Zie5
sTfuGRcXMoXsYOz41JBBhTYbalOzuIdJJd9Qs6fP2sVDy7tbxnWJSO4HgaFLBcb7Pj/LIFR8YJgz
sPfeiaKsqEhrt3MtubD6zEJw/bbKYPQWksrJnYUDaAUu+S6tgknXxIFQubpNMF+yiSg+g97MwFwx
3lN/GSNw9gjhR3FdleBKRP+kMlntY4yc9pg0iVAhggIaO53pJRYfWeUMiNrlw2La5MR5qUXql1st
lzBO904f3ERYHk4H9KP1Ts43F1nId4EknQT93/U2ZAf9VKkHtY5s0EUFaIbDurPNAIPS13BUeZP4
5q1D/oyuwd0nPh8bUvVuxSj6WXytmJ4K/cvJvCp5DeCCs02BL5e6PJMgCSq/nWAidweBnvbi7Wip
2ILriOiX/glkqa0XIfBXhdnajfjOZTHg7hvadpjp2NlkoKjBk3FU5DWTwJkSk1SnJ6U5xm/bIEsr
Yz9awX7Gu0xhuNupBvymJy2vmQ3PQ7q1jhhLygkTTK8+QBozWDbZliLTGzYwwNSewd61pXbrGnwd
l8QJLT+bQjtoefwzdzMxiEYTfvOm7WqYYY7cj41QMqR+X9bAcG1CTFsTXsEFVWNlxgQlW+Tknqbu
aMsruXPnPGnCztavIxX8ZzJGllgvrfHAMFxxhyc9eH/zlA7LTLWq+6ebQ3psRMl9Qiz0YYIS5RNk
ya3eqWQhgSmqJ/H0CrXksBb8wJpAdXzXXEpdySYwXEWR2aX6ol3poOv65i4Bek3Sv4EMS2muHqhA
DukiMBDd7u5/9D0aLEtGQnYahhwsrBPUteKqjvUa8fdNWA2GGwvpTzKDBaZ8vUZE5agLK1PJ0JY/
4vyzCX/G0ig5beGagAg7OAg3bT824rmBzjjbukeLNqaWceROSHr9McFd264rZ/Offrxv7sEu8l+J
0FcAKro8TIhT2SVYIxjmxGToEvBqbg1VJwqSOEaEpNIWHWRWioB6EpwzOWqE2mPoHjKttifdMUDg
uhH5F3BgEggJkh/+uOUNza87kygPplhqIasmTsqSEzGLYWxuLo0YE5JsGNblpLNfH1Jbi3sDb5Sk
6TdAXHHNCHfPEwYas8lX0g7nkDAAJuSt9R4HzlnVRfcmm9USHxy+1oJWVOl/Yi99pg09OMo3PkzQ
6cNs/Rvsx2xvePD1RirTrGvLSkNzVTxT2XX24Tq8Z4lFsJQ4MsFAD2IrYJqx+uhK7AT8YeFaSe+v
woOxxbDLCd4kLP4q1F7I3OBXdYqfd0dzVDJAY3vtw6UJ51U/5xesFC5tNHLGNFsXmrUr8oBhIQuj
VpdwW5H86sVDRuwnidHzbcJOfTKF4IqxosDVstq/doyMl8ZDvuFi7PldX15KvBjpkQmBwMduz3Yi
Lk7tqJ5yYRsAOaarSwVp7vXbxcT/RrJTubx1S/x9XN4ava7NU/kKY7qXCx7yPz50323u5UzPLxET
KMPHeymCPnUP5SbgLy6kZafUFbEjMzXisovDtlrVtCK5UGRYDKoBhawmvFlznuF9OuBXM1/pn1sv
JmQ8y4g0zv1BznnV39zIVoZ6Z2Ru3jAEPpRIY7WjPIF9HXsxNq3ZtqHbmMLVdFxNYWE4sgNoivbu
Kh9JD11coYxwLV/hNCPHNyZoqs2IF8PmEEF9zFDHv13TeLiT61Iox7rltj+UIQXRnVL/NyYzskXo
vlw8AmSbkreVon9rGQ06zBJQ7+ZnAyY/WTDXi5KLEpXZmmD0CVcvDW0Tn/fH/ysCeLMKYu8E6tZs
pjw0Jo5VLp56JEBIVCFMBWWZBaYP4pmH+BUGObAp1eV3UumhsEc8ypoYpFNEOzxnNbE3hHqaf9Ea
msc2CD3tRh0FfSbo0Vso1whAXKiviajioMWEb2iI1d7yLl+opHNJNtEIlHvJrH2SAqdvyEe5Tw8O
YhVhG2Jg/eAPuheffUM8Vzfjkzy1c5bTIvVakNuKWOpZVSpNE6QGccNWZIbEN9C1lWCk8kInaL6w
UvDx0TL0EhxkDl2iGAicRgg+XZtXXYHIfafbPLaca6r8n7ojG3bdA22LVMTgc/6R7huRfq3l5r3i
x8By29VYZj7q8MJhZ23WApiXjbyqxr+McWmG+xFI7lz66+9TZFYy8Oh++zmp2mW9GnTn2/g0mqaa
fuaq/jUUKfmf+vETqd+mK2YTKH0jR0poLaRYOydiGJoRE3BEOCzUiZnUYxIJ0jhTM8pLNI/gOLZ6
Tv81hLGoRtv3cFKsigI4jkNOrZJAe7uEl/JHWQUI1b4Wq23QKJk7xURupZkc0XHLdLLBtPOm3b0t
rxBmiThaB6+FApQYVhdxciIpxYmnrreshTWLDFJZfHAmsuvbKBYcx57iv32PB91q3ZuzyPS4CUJW
CrnD0qHJo056AJfrHdp/eIX4ypDG7Y1S4sa2Uj+FmIHFcfzJqUSfL+pY5TImgKcp097bUvA+qCoJ
sctSJ8ByhkpOnjBdh6EcvUKpA7r+0hPbgReo0KIofdt6TpvB7+dMn2ZWMUKbb/ZDGNuGmrhcBGER
GLBnzIuSTZO1hbd5yYbW8MbSC+sI98gd4qNs/hpGJSiHVs1YYizgLnCgYH6WXOHEnvgJH0csnm8y
lLMbmnA/M62tQaNpKEOXVqxGo8SIZAVOnY4tyoQPcFiNIGlZwzjQsqMhxGiIZxhhObQ3yeqx3p6T
rb1KxX30SsZeNx+H9n+8qzMj7CN+A8bbju5NPX5xl1dzh7Is27I7/ZwiN2Dh3D5UmP8pl7Mtax9w
6612CrS0VnQNw5OGBBZE6VFI6DkKYDh1fNE0437VOirgMZ7E1g9uBAgPWZsk9My6+dBGmuM47aDQ
CMukJ6sAJvQP7GIrSkJn1n9r9jJ2uPngH2i/ndETfCXWChMk65AkmbRduB/a2SJfShG4SQknJrr/
WlmNJkmRfAdpKyEjW5W4s8W3VsxxH0lJZVFYpHn9dmRrzOJ1xQOTXeAx9lmldaGViM/4ZSPkE/c2
JFAX/jYCp7Jlg5mO/DVsWdd/DOVSEMzPohaQ3lv3yuxe7hgf9RnH4SGN5DHOlYcfnOV2e43LFJTB
XGwRyl14avvU5CT5ktiGG3Y4JFysWhjr8s/Co2lbUg3loEbfxefl8SP14HJqmsMivTnL29tiL73L
D7YG3nFiya20shYcHO66KPA6lyf+GA4iGbtiVfRH2RjDQmUYvVS0qiG9t9BnwScE1Ttputw9YuSk
ThE6QM8i3PVf29/XVBSkZvNkPOpXs0NwCsvufdgysCM6w0S+Dp/896eTnYvxoj5ZzdrO8j/gtW0M
WWwByBMyaSc+/mig/1ylXjombYe2q0ezI4vp6e+JGnIjpMLVGq/17DpYcUrGG5RqGyHzjbyyhy+U
n4yQ+7YPn4eyJPfj+D936mjrj8fzK/jPmFxCOCoDxZz9Fl6xve/8CK6IhTnpXy4RbXQY5C/iQD3S
UdtIgISgTX52zyeMtmTQ57bvgZbfQwwgJL0EU6IDR1caLxfoA2X0VfCO7wJ2qyrkXzshxOZO215i
aQmAknSPAMX+H2F9lpY8KOl5xN9Byqaf0/fXLppeuYYXZMNl4WQ3F4D9OFPUciiUjTBoOsbtHeEm
+IJxBXUUQNKXvemnFmVGQ6e09q/3aRvtCnpxcv91gxEc04nDazvE7WFabzaszqj6wrGyaGGgCZfM
iJ6ZhzaDH7lt4i9amq4dCh2AczuabosT9FNNfc4twe0+SvPRrNx+bUJiySXnAuTixlRvZZIa1R3I
tjFuMbNBh1YpeyF+wsqyyCtlmX5WVpodgUx3X+mhmyMeNgDIaD2MFbx1Eh4UON8Zk9MvMwrJ4tNQ
EUsnTrZQ/kNNHowSyln5MXo93p4kaPy4hC9j0zGtHeIJJUmuvobT568YQ6//4n1p99Mgq/54CoKi
BUc4PrkH63YeuDdwzzQJWRVdwO9ZYoWsjt52IR0az2Ea2nxnliJJlCN6t8hbASlQepVSfC5BtYYb
+BwsYzNYlBbnNl72hfU6eSgcrhhqRm+ZMm4fOfE70XFF6gYMM1ORngJWsTGhcz+gV1mKnqKqYVYj
9kvMfQY0NJhyV2uaVVH+1YTbqo2hg7oXN3DkzQLyMqHyk5N1aiXvrYKG7v6yAdgk9hhggCaF800/
5uuTcWWAAJFtE6E/GxjmsT9Zvigd837EMDk2NKvojZz5xo4Pnl3fPKC04zeIQ/uUJ9K6C+cfHlOK
SEfe61bW1qa6Mu4grZP/vaeC75M2ShnSXqu1IQUz6yG+e//8zJnCn/2Do9D8hM0okbvKBLDWQp2P
Wb8xKkcdPp+amym6yOLhcATf8iV1IAdDaRNVYxojiAie2NkOMbG3l6DNomjuT1O5+02NYOytE6Rq
BYmrz97Am7f6w6N6p/6BGP+x4nJjECXyOsPxpdAMoCSkyw4WZAV4NFIADd9sjCcS0I33FO1ja+Zb
pjLct+ETbryrzVL6W5nsYReQVOHsNlu6ag66nlhYERaJ85vVjwgQljMJSxKl5rComiaRlM9barvz
KdLEw/hrcwAg+FgyynEJI8wvhoZomtVLyuEj9i0iGuZIcT0Pue4ivFLbaAfMCFhdNPbZMNRnI5E5
DsTE1DwSYd3n2kAZ5zkCt7qv9cUv6Kes5RGKhgTsQ5PeFckdqj8QLhKSX8/K1/6latEYaIBJz1Je
LKVqHQv7mH+0Y8i/ir5Hq7sj8MBuHTluslLd9kEsWLxyy4745z5KdtwXVRGv1L278CoXTYCM3JlL
ObRQILn9OwDMRHwgVgM8VG3In54xhmt9qAjD+Q0NnHzilXJRvIUREwQc29FtyxdnOITr520nxEgg
l4/R2O7zLZ5gB17erZEmGGZ/kTjv5jcyKuc5SETuzwvHRDo/O7OR2HZgrE+MU/C28GUiEt2VLHVv
vOipIlo7BB811+LKpDWb4iGsudUFUyypzodyzetolT+spzFTHuMNDLUjYRaRxM4744gIryDy+heZ
Bc+DtUce13djCyxIxcL2NqrVJqztJC73wxcVvgEQde8S3hgt4px8lS2e2Q22s9d+5FTKpda+hbKz
2kIlDeK6UUeohcfV+MjZ8WVM7hhTZzs7w2hihBDjNEeEQoikCoyIFXbCYEnvMwhkItmkX+uoR9gR
o6tRX8u7PiKejchsM5dmad1J0qpkJmiDDLVnL67wNE4WsrZcz74nbylth1kzwmdIP08qFfOyOyh/
a4yqexwaM40ZMARc5KP8Uskh8mpz2gxQxp2eXAH2w994DNxcPZq7mx88aDS7oUxvgnLrMv35hnax
0+ShG2r2cCETQvflDLcqWUqY1IS0wOxUs+yCA8J7a9sIOUYfbPyGJ5S0Hv6Mq+Rm/I+TnM7dhhzC
RphWTa2Por6HyyR9dqPStrUen7JD3JCTRGvfawR5NDI62J0VFeLmFpbo0n1tYmh9dZI8JsZD6kpZ
GPjIo/aMpD2ciyrpW1mwrErZ/63LRqEjPcROXhGYEJvCmjbOxrsvqH9bcL/p0mA56O+sz8RuOAhU
BWazDvWlm9dhCQfm2s+qkUeaMObhAPJgYmSIFDPdkfvYXJIz07fu36cxEaUTlSCiCspjyER8MDvl
1gtohB+ajuvUPI1+OL8t0NqOelE1brN4OcZYn9NkypAGXN1DTTyiHBqmi90nUhIessiRY2qwCPNt
u9VmEVM0PkFTf1ephoLIUzlpuPqiohxrQIZrEPsZVZEcdlROCYlS/mu+Xw6NSZ2nZ7Om2osUuv4J
qzD0xaKhLcypByPu4SL/bkUNEVn0wOePt0HeT8RhJxouPqqga27rY3v/RIvrPjsTCYYsLu1vGHDq
vjS5SoQqOLYWlJeHrMUfKBIs+nxYHSTh8yO/83Q4litT+hEDc7mznLgVlDHnUPEkl3ZSIl1HYhjx
KS5JjIIZCpDmeGvhEXiPVPcHyBcY4Vj+ZgtVsnWi50SM3IsAIAgIoqAEGoE29VHfqvVHdlTIIMKh
rJNpNUxHO8ZpsBA/S8QIirJNF+cnM5cWx7XwLcq9S/kcgO4nA3yARnLGTaVNNhck9K2FYFMDaYNc
OM/TXO6H3aV87ZGuAzL4QfBSHKXkHXtP9OBfMH8XlexUBy6ZoeaJxtCBhHgwd5CIyQdEcjC0LHE9
GNY9qnq19eigDo4tdmAnlEnl8pYaDj3qfgSQgy2X0dKMDcpTp6Vt7+OcpeU/qvLO2GG8Te6L3ePO
tvdUCCCZ3JCBfFGYYx9zl6rNAT/0rCRki4VaaHl3FotucGnrhF/U2W1WIK96w/W4RMJxVjKasyRn
UD0pgGSc9UcEaoisRoIhyEm+B/fMNPCtM4m5hxUeuEpVwpciEzRO+Ps1JRMZPXl5TEYdXuNJqImQ
Fp5JhjfGvJskrOnaKM0nb81eLAA8y0zoVqRgez8zxL0ZcyqMLo3qpXox/KLn1yq6J9/ytdGfDjZw
CzN3AyPvjgy0P/I69JGqR8FzEjzok49ZQBiQx+uNXRLnnkUjFCQTRr99dl8qQ+57g6wNNuwln7bf
9MbsyQd1VoThuhqLh7ZIe6RNZAUO1pwvCSK6l6F0MhZtdMjf/46Qjqpt9eI4o6YoD4imVMV58i0q
nfxKJj1Ft8zU0eIjiTh5BGsRV/wk0yMZluQYdyOlAMH/agpzlhxHWvnyr7DvDVmDW86+cbRhVzNK
RfjJYf35EZY31xcnTMtYvHkH+/ofPL5FpHdy3Qpfmft+qB/1chsoKB6CXo87MxB3p7/y7rRxnjcd
YYyqrz5uEoZh6a2KCfsGDerWL5it0DsSKxgn2hX5OQo8/w4NtWoB2TmJ0yOdZXtGE0OA/g1csBhM
LfQiO8aRGWQHxphEEjcJwwvXLYmJhsfdPxHLtc2BASQF969Y6JNlr2AMx1js9hZja4YJLCX0sCkJ
sX+MaiGm2CgHxsKcNyyGG5AMHdcyNCZzX6lRil2gRmHN3l6EXaA1q9wBmLgU64kBWszXiPtH2fXV
MF9NGtmxd3vig6XhvwnoBq4ve8WQprkvFMwTYVdSYo433Dm9ZOnH2VBUbvTRIk00dyYRbtD2hq5q
WytCi0ZZHJtGRMms7MtM7ZCBuMuujlcodf0PUTrk5aKZZJqnsmb2WLTcYBNneOoSEwWtX8lX4dpA
2VsN7J73CABHzNxS0hRnLEQ7VS3ytfnuf+c/x0EdM9iTos2ZbhQI08HF3rzvc5nHE1IwcATfxjpe
0mvv1j8siUJOqMgH1cEPHZF9Wl1NhNibM/0fcSHZZPXLd3nXJ9IdoAZ/6Oa5JqbNz1f7G40jiB2x
720504BU21836uOPyq0Jyob8z2Y9hRpxl9kxMtYvaMqpSffBW6041GICPTjkp8OqGCII9JN6KZt0
vOMFyYen0gXABu7ZFElm6uUeeRHbzpOzZenOSH/mJ5kOXM/H+5fn+BSLhaN71HTjwLE3P+1WdgKU
GLsqJpVQh4AoUwU9E2v65QTKKnIV0hRKrud6PmYnFFCJzPJ1r/mAQa+as2Om0U/ZEBYWOvH/wmHl
zAEVtGY3rbeDR44tWmqWqF5iRvf8vAa9Kb/St0rA++A+k3Ga5/v+dMWcKkNsWRmGMHEo6nEEUWMJ
j3B0M2rwCB2gqhvP3+gND5Ace1q7ntR4R43omLTG4ziNGkUo+ioapKLQH4qiVq/efHEUjSmwcovx
pqf1sl/pmhdh22vX2BrrbAOxWd8sJ5tEKg2g2d6vS4rqXlhsKmJI+qhz2vTFfjbSt5hot5vTD6oP
F0KUqr66bVDVXSoCfK7PixC3W68OngxT51TisEe11pdDkIgucvqk7R8sw1dfVX0MmO9sBGL69+Dw
UpfH5eiapcsRbHpldANmgPmqv0waSbq3slY/ZG93vLjxlIyZMTBwLo4M5Sy1Vbnt2MsszuNxvR5o
aHTE6zDtXV+iAVEGsQ5woeOi4Ou11cUbKK6UfEa4ozDPPN9tj/YgZqeCoQvF2gZ3XFfbSN87Kdli
GeYe/dC+8XvzyWfBy4anBihUqwuQrVnoHQDyJKcevEy2P0pci4wV+Nz+2vQXsWAop/7Hx3WzipbY
zngPXMowqQ/69ioknDmIr6FtWneyReHmzwnuBJZglPiCxNZktQFUloMvb6qbmQo2MZDrszT6uX3Z
EO5xucZmx8ycZ75IDGDZPNRIptzav+I5f/TC7Q7/FWYEsckfq6Nb7DxggL3veFRbp2MK2lz8EHKl
nVs5tbZNPyWgKHCuJrW6YxzjFMc2cAbkZOdaz+hp+1baIGgcxsV8uZgxhA9QrFE4xR1N7mzH+bbj
74SRwywlK0e41juvwdH8lEAGPKKi6GQ9V4CcnY/8p+ORtCdbnv+7e+bAkQd9h/WIc1ytjhfhC/uh
JhVu1iWou+dWATskvaJgz7ELmd40L6yw3+5b/bL5Gz3GczXxkL5Y3WMYVi90Zx6U637SLtZPnmMG
VAsJL7WCTbo2oYwLYjvfBLWrRhk2zccEUSuqK9/XJthDe31EG1V3UmLSMghzZwj/egSFET0iJW2F
NW5LuqZdNC4EPqXTjUYHbL7gJ8bwrB4s74dwZP9uz9IEHvawYedbIBoaxWc2tKRDgAYc8UrBJFon
y1RDAdmHEAgS8HpecF0PXspwbgk14ILNUfKkfl9LvkONECeZo1NZFlLomP77NTCtI8CluYN6Caeh
z31MMKx27M2qXYxwSPGpTIS8EolYXC/u4/fDnG8Jpe0taz/aP8by9EQNrPP4+1EpPjQLQmwPLdhb
XsMF3OHyMqTRjGYK2hzlKyB5l+Puq9932TpUdID89WpxocDaSoVEynd2J73n4t+tPkKbvhsCPWyz
GNC5EjaGYClMzbesy2sm1VGo0TMrxvc9JCoJ6Z9MclArh/MZbHGl2ABrCorA0BSD6gmoYW7AFbOK
22qY38HsPNPweCjVs7F4jtksZ4l3fIulCyqJEpXlZc9GIxT2DYATGQwB/0Wn+MeteahNrJ/XM0dQ
1+CqycV5Y7I3haHTs2ChP4oQzJyqA942WKHXhox1+DV3LELudF387mlpNyrGYhUEaQIqnPyqGQ2D
feDhc+UAjLc1LhHc7HBVstg6TM+T0/11YTFw8vAsBdo//qx47M/lW4L7ohpbgghkfBfY0nlvzn9C
MPX83i/IYQ6wCZsiG1TKnw+CmQMslLBqGKRemWeSNmYnSqk0H/GiZg4kNQW6cw34mHFaN2/kpVPu
cgZaPEiT2KTqn3aWJsFom0H0BzpbPm0J2XkadFAhxHRPOIVvshbftZljyuESSb8Yq3k4hZZiEr5r
7yiieeJKDCW2ggnfcEbiQCNKjh6QA7WJVFH5fUSS/q5FnKOdA082eBE+MDgVIptAfH5rCKCkjvp3
2QZwwRQVFk+Ga6YykgeAvPxnsgyepxTvW9iXzkM9eE/xw+8wY8Pkb2Xm3sFqGZFmYCF5IDlKgVnb
Qzf2tug/A5AA9PYvD6Oe/UKzCc2q5dz4/5juyvBj36B0OZq8QeK5qqd8HY0QuIJyNnWvQEnk3fvT
m0evV4gIPcCx9L9HDiaEq6KqgREs8m2OZgYwhwZkIxBn0cMQMXEd1qS1TMrcFJqE0dYXko3Vt3Fb
qQyeFu+G8+T6vterBF/a4lu3zG4+ukZIPO1QomOntw+6m9cTDe9kVRoVmBpos4/n0UwIdLXurg0h
6y37YpkgzFYz2y80T5O9BVjTNh011qBQL8fxoec2fm3GxA3qLkcxuFAIl7hKw85JXt2iGRHDX+0e
XdVitLCFtR0UDu0iqs1hSlKd8QafFrr+EKnYQVVDtmA7H6KU4bl3+U9B873S+aobDmk0S2xKYXKP
xQFh3ouGqsqCWM5p31vSXXowsV2ZGZjztO4VjhRdtrDdbcbkRDGbreSSVGG9vWwkKsLQzA8jhMeO
AXjz0fDSYZvVRhv+vHUd8fbs22yOTKO+91LTZIPnSz4R7/jVwCDXDRKX4eNzPVhtvDhHxGAf9GEw
XgffTpVqeoVpEsJoXCioN39sIYx+aH328l+D73s7UpwYXRSUKy7N2u5FpHr4rDSla0m/oWEyJgoz
GVT9FLiO//NjHLLltyoXrpz9Aymc8iSqUBgMv+Tj+on1QF3+tIEJZYwFhae8EoMeA/x1xYmzqVbW
Keo5zpvsIz6e0un2lixzuc/iANJq8vrZFPz1Ti9ufvO/Y7ta1FuzQl9LWc41/PZYF7G9NA65olIG
Ha2lCVnfQGUzEIA7HUirYVE5V1TNrY4KsgDGHiQ/0Cj3+WXNmbpa/RVHM+WjbKrDohCIsSxgkqTM
YqHFeE02vh2XzyBqmwZfGiyUmKPt7Spuom659CuSm2ehYKfqIBbdfY/TrQiIdY4rhcED7lLR/xJ7
oLFeu1W7rmFwnMArkSs/XkSZq+uAlDZVUfdEDKjDwd17oExdRiIjwMvyUVAm+vRovkYTvRW+szLV
nXtoUbeOSYDw65kRGJHtCEMmXgEZ6BRUhMAtfwaWBjcVBmxQuoNzT/fHCcsiEMQrKDNYWhtVlX9K
U2EJjXR+HSp5dVws56VsJfWDBra7OnjBJ5XZ5Okht+wVQvV0yFGRNYWFqAidMt/rgCkOSr8rliyF
ndcwQ5FxnZGdAzw8Z70nFJIyfUHDxgTZ/kD56slAP0ny9ezqRd8L1shKcuoRkVpQ6m7twJBfpc/W
3MEDxMGbUWnFGfr8ki3/GnViHs1fk8pBLrv3IQpDfvuiFX4Wj60BjSjEQNdeNBN/N1sR3B2DCYf/
+ABmIYk0/4MAYKVzyArJeoIRoVf4b7TsPN3xrsm2yyqw68YIAZzyOR4f7gbYiIWafCMua3kVQjiA
pt29337Ujhw2jcy2YmyVOZZ+QxazbLVlpWkvabEjF/kUFBdjI0AMdL2Z25/xB3Wk1WstYTT5iFp9
9oJyGFKc3FW+T9HmMTwmzkuKLoE2FQMJM6nU4eykemWeYjV0erGLw3zP6k93Es4Zz5pXMESmRxxO
J6fOuawTvjX1Y/0RyGxtXW9I1dByfKcRpzbiUxxJtIIhPyI1gLVgOEunzn/y0qQeRZolkm6V4IMf
O0I97RTpUsqtkUo/YYVDsDEzRRchsOIXn7SaMagjTGyrImAADdMByGpgKEZsEP2gEJxxpYxdpPmT
xblZvre1rA3Hg/KRu7hMT8o7lbrZeePOERnqkPPT6LhsvVn/6vj6rTsditTlxhfNv/n5Nph8m5KV
70SyQYF/gqmFaw2/kT4jvuu+tDwaKxuNIaQz28qMMZ/A2kS78D4OlietXzjIiQolkXvcl5oRKq6Z
dEw9rtUoVVOWJ2bj6heEOVdswU/GAlvbnjk2Fe+qY/3IS871Eo/jOZjcseVbEJ7BKIwvo31BcTSf
KhUOK7Vtdr/Kg3a336yvzdKovn9IVER8uFFLcBovJHFrke42GdLDyBY+0jt6Yr39KMZqEIxq7Z7h
f3AcOJAfS8zgOopycJ0pLRq7rDTbQkzeSMEP5JmBDtG9gw/Sjygn7NbQTz1mbEptYlblfFFpI13r
KQQC1NZBPTvbJkoGixJow4Nea8uh5+e/8oUDSHJSe80OMP5WXu+6mmnyx7mzfb/F+Vzg5aeLAjxs
MmdwawGAqiiLjZmC4ViJWnjwh9Htto/lbPtjcaD0Wm1JR9/S/ha0pk3uxFI+Ayagzm4sw0qao+1R
ajrKqsMW6LyJpBlHew+CF55r0ZRvENRlm3h8SZCLIy2ZImCPKgeYUfUrf3MYhjuUbBOsivBSb0tY
0VsKfbldiIpYfHEAU/fzrfyDyhmqYEgwfEu2Y4+UnshYlbXXwplu4saylFRwD4QHR+COKygLvV7x
MjfNOPrbpHrOBbHuCh6RLd9dArD2Sack9F/4tS04d1gp6X8juiEM4UXSJiUELhGbV3wOAXEVKELg
VQi66yKeoAUJQ+SZSuKMroemGRw6opGHkMhHcsP474RUZrXyBAnNpy55sgSJR6f4PYKHRt2Vquut
nJKAaYv/zIxCjhxqccTxzng6VLeiXv/oSOKRLKa1j0T6p0XQf03KMqIJsZkg02PZTOh3sVPPb9zt
25gfW44CQQJ/oShvPI19TWPEwHK5uzboVTX0ugZqtI9hpm24lH/5zZ/7x+l6fyKCuwaxdBHo8uQN
SEpA1DIVu4LLRHsjF8SiROccFHJJ+kAUqjsIuDYSr2nTKSTNANmcy4rJK/Q3bd18fXFYfkaoUHf/
4/xNWEtOW3a78qYQ6xDVf9ZBfOo1+5eMqikUL01VxlA+i7+ATSVn1q8NMEt5y+iOKKmgetcjuZ4M
+ZVmTkJFnhm/Jnoda6B9Y6qOWmhgA9iNbobUIOirff1jQp/AAbmmQ0chJsvUwNXuvBPpGq2+ZlJR
JnXQ44lmxlT55f4d/grUpcK99e0GmUcKNgDAu80flDQ5URU16AfCwQBbpmB6SPhjubCoYep8oPEs
G+Te7M10I2bp7cYPBcpI6RxManXWJbgAREEK/cp0lu4n7Jt0T7RLjpAD9H67KIiBPaRksA0C+/LD
pM9+zNPVlzQbNR7d1vH96AngMTuxnU2nGh1MiZSl6Y2+lw+rOfNSJ+2Vm0ncDezkn6w/uUpQjcjX
lSQDVMwfo+jNki9onO9yu5vexsK3Wb3COUCKTXIZny2PInQ/M9YDxu89g3+GgCfybat4BQcUGpZV
8lItG04Gg5Bbu3bUFoLlrZBcWg8mUKfXHvMz3vAumS6/V6kJq66I2T9dD6vVyrzRIAztk670h3HH
d6wdecKlF8cImLMNYi/zyXf9Gg0MKLgRcIGaouYRPM9fOsOI4hvOzVzmFfrRnLoSPVcJtr7aG7c8
3XQUCnlV29VzSuC4m2rJDWzb1GMvxpVLEJJlONaXR2UwJ7XA97XQf6RPuuj6UkSOKw+fVFtFHuLo
XCd1ThXgVqFjc/ov6dhYQt+kVQAAebkEcsSs7E6mrTyWut0MOLWMIXZAFrGHHRNdZsxhcoiviX3I
qGo0ZNBkeJcInzRWy/aCBK79fngsM0HnQ6KszRaF0bAFGaO6HYSvogveD7l79GxXW/zTOiDj3I/Q
SIZi9VvMpaMRm18xIKV/SdsfZqMh5+tX0qolArty7Bp/iPrJj3wLa7EWBr4jOrEQ2hHYjKqAYqf1
CuTfiiIoHf84GbndfIAPkOmTgPoZ11BDYF+w5O8xAnonKl9Yf/PiAQz2mPh4+y4hL3mtkBANTRMF
Pl7XrJDZSQFo6NDBVUCocF2OTRR7oKaT4vAU29lFlaxdWxO9QEpLQIsYjo1ZvPpgMNRBwu4LrbbU
LdffeNhnwv3Og99fZSnHKerT0FLAe57TsOow9sMLhH98zMIKmkM6n50KHcNHNI43O3tYZDA9W6i7
kvOkPzn3H5mxHTjfq4PjvchTLEBAok4cNrKTMvxKrzeGyoGzGp78Uiyalgk08Mlto+PwatET6y/5
8tUgZQ/faStwhW5sG86S1qjURPtF9HDKXhcF7FXP8T+T0B2MKBeKi1f4E9D9YXI0uTuojl8WSBmm
Jw9hf5mNYJ5K0XF/0rpSQK603xo+1rcjXrYK8u6jjrY698F3KFIU7Onm6dnpES4uI2bJt/a6Wxp0
6tTlMonz8HINP1BS6F/lr9X6VmCCfsSMg4x1qcH6wXUmHb3EKNtMiXxTFaBl00Cw+XS738tIHwVe
m7FJbizR9Nma2rbluB7wmSY5Y1ZNz0Ymf6Fzrv1kOO1pygkzQ1JOQ9EwJCkY+1t0epcHmXlH4kGT
g/s8g/hGCjoi6kiSbmQ/AOIJ3o/4krlM4CyhRCEavNi9jsnXPV45z9x2ooMoDBjMHRzBdVICK1Kc
WgYHkJ5mPLOfCs4qa5AMqTeaEueT71H7gYCgj4KdsiHNM3zJzlTvq3OHhGkr0nUnj1R/Ui0I+2y0
stb5gtoYw1yHgYPLwJYyN8PmA0juTpqEDa0wnZng/bJ3PchZRr3oclPD+dzc5TflW64PeFaIeMbw
JEhUTrBT2gPPeb8wTP9lHqP1jwGrQYvHBCUznNecULAkAv7BdQJOwUa6qgtI7mWtjfjY6mRHkjwT
AMzw1KjI/kYLoC8YV0ThdbDvHt8b9iXv0+fv8kroOxH/z9xnMaJ22zA0JWHCWLHmnL479YJBgA9E
URmQ+LYe6sj9KS1jU9PwYpOV5CXS7ic6HhfctusBBj/HAc69+sFUs77IGNFD/AZrR1gPq0CO053u
0dAOXIx2etllH3GBf4O8ZYm62NBiSyicW5cRkI2uxcH1G/N+NydEa6I7mglEmR9G3I3oiUKp3jJo
+wftHv2li9Ll6P++L5pzcD0A6iet9uKUA4uw0XFhj5zH/DDHuNP8erCIhVDHQfyC0uPCRFsHHYMP
5ak/GzUKq6dzUTb96E7UilqvX9T+2b4w4rO+h1Ip/YM4TZ90cyG2Jz1okFqoyvp6lltgWxJHQfpT
PwnJWUWlXAZZjeoAzqxEVljRbIbhIeRd6cKFigw4gWpbkAdh3sk8QGkFQtEg1H5sxetAeXlRLzaM
MQHgfUYAM9fVda0nEuuwbfSL11iX3o91HT/VSwHF51njQn1fsTilQqLIBCTU2h25KdmtwqK6btrh
2xhTWuzZ4VQ4dc72p2LcgE/xJ4zu00XBjXm8h6Gb4UdCNxApIJhmP9G8++LxU2PTCIft5nFXVxBL
4peCEBKFJP/a4d+GnRNIDv6ms0PDauSaQqlFvKJcM0V0XQXgdwuk3tnHmrV2RO3R6vvi0BP7SIpZ
QWIRjJ8N9Sd5ZiRG7znRR5NCzsXTRYlCf55mqK+rZtbD/TO/Z7m81foOC0kje97JiKi2MqohJbgW
m8nxrIIOOkis3hKxv1HLx6O+KoPneoX3K5lOQ2+IWV6R87ANZSxS0zzd1BhQPtATcF2TWLy8rQpl
GUVNUtlgT2ucOUJnZ3axlxxvkYed7k6dBiB/LkK1gO6pYN/EQKdG5Ny/52rK4MZwcf4pWkwxdU+i
1RrFJYbjCUJJg5Zb76pkLC1wIWNdIcKtPrX/esL1NV8k6ddlwk6Vdtn/a6tCOzRl9BnhD7mXaPzO
KnJLpXzuGv7lrgaHLB30g10PrBDCiPUC7ZHhz/gehBwhRFLNWuQmRo47KnEpIExWoL/tV5WkHf5Q
f11AlEeFp81mfQAQFhDDh5Je8Ag2nQGPa5W3zt4a5Zj45noHu+vaK6r/+d+YYYgntlVkSXWCAIBN
iMcwRpA9dxniIXVvrILsfK59vJjvixso5EUZIzByUDwU/z6A8bamBgPb+RXez9LZvAn/3DsMsb51
fL+lfaiT7sNO+unf5PxZgm3KuzhbUjZipCT7XZV70Fuook5EZlZFVZCCy8jzupp5Xv7WLkl+3M06
TaBXz8e2A/FgSAMImdLqKyIwl9Jaa5jEWZ+euRM7TZ/vHy4MwcZbI9iSRF7QF2L1OFpfl8c7go5B
fCHR7dXug8Yd75cGZ8DgpKhKUZP7tUFDu6/ynKoah5it1zWCPDyV+Hlr5BziKX9out/EXXk6kHDH
iXSL6VYyhcd1VePAZUtsU7AF6rco1Xy7C2ZEgvPRohkdvWeA+PGTaW61Rmnaf/izlb0zGJB2NxQu
fUL43Sm/P2xQybcJysb5MOFU2MuwafYOyp+m77bq7TriakPZRNlzQv4ozScSiZL6NDGZ5QYBNtI5
0oyTeph3zAxAx0W3YK1awKV+Z3YD7X2ZUnFNjj1aKjFGkbE0Hdy/po6aqrP6NBR69Uuz2fVeSNjC
zrF3b5lj1TJbp4Pshca48zAlCZJsHZScG+JColUooat9XV3oHRWYTGmjea9uI+TOwKBWve57/mjP
xedp88Fd8yHOQeYjG1901RWVdNSWbS3nGDHpoQT2zFelE/jOypL8/r2i1DQXRUAycp+NRL6O3zf4
SkB1gjqCIDVXJRxb44+q8BysnQN3a4/418uvnxLgPgGZkGQu9gaEOhdYzwNnX3v+9ZDehzO+4+Xe
4PqxzUNImI6N3IGaob9zTDyvfUQlK0udW9Qaq1F2DmLAnPVtG/djuQj5c/Ik73ApJ6V/rwWV1QmJ
56RZlwXCIFGRTYsAr6KUm3xIKgaOZkT7vf3+JM+QH/mdlRs5K8MdBn6ND7vfcPhZUxvmNMY1EaCd
1fGPaGa1wMnsoEzUywnP6eXi1XIm++N8byJfeTX4Lvnaef41wChTlXzpVuE+BF3ph2IVbZiwf1PV
3+4+EwJUNYRCAmGrbUGPZ7xjsXqrTTNJJijWui7YpaT8of5IyJpkJfNJyutbilHBALFjVNvua1dX
UE4fvxVBk2jB2nrrEXYCBxWH5ib3XQhmDrbHqn1ycBR8MLhNgrSYpTuLH/UcxTBTMob90rJ0nanr
AUmuYCL92M+YYRsU/KExcl3llAmn4si7+Eps7jNKrRRggT6/Az9JQOwH/yD/1vFkHuZz0gyTknSw
pUBVlu8riz4bX153B/PbGFH0eu0kAGtO9BezFSrhxqfX+BIhoZEw9FQCU+rMKGYrBoCfCIKFVc5M
cMBza7+M/2chYsfVzdJ4KADW/qf7aeQltbMQnnLeSn8hP0z487uXqraemaxbwIxTRHOVKQEx5ZuP
HYJK/zL8qSrCHOMCDnZFztu9aes7PzE7eZFMepKb8B0+hVTFYaFXJtMjWcS0kdPE5v3VE/U7B3X9
+obF/QleKr8wZ2LvhvMG/S25xghQmD7sF+5rKOxOrILgZ1hWGa8jCuAT+6cFCGxgPgYvii2V5KL5
8Nw9H3TenYSmESvJV9NGnR/3oeaooPIExoKZKOymKkXRmp6s+/oP8w9zhC0UCkoefE1zF84OPYLG
a1zbwpYfJls8BxyLclNCi10WxsEWmN3j4uSomD+GhC7z5zfuQLZqiVqcX9vOPepVsGw7R0KS5oyA
9JFzYVgCOzL3tS8ckFKkKW4++f7WXmYJXC5V/4Ej9iBmaJehSGAC8GibEA5AwsyFgLJmrUHMzWkq
NjsdwAZfIX5n3XjmjBD0hfu4owwWRz4bNSVPFKxuKtVzt25OoTMHynCil5ZgH10MY2Vy4BStsCFl
A6jpTGiSrADpSywsVsZ9YPU0gnnnfS9zO040YFNHYYGtdUIqJa4Uo6JM8RfvBj5KD0pEYhm31Oft
jEDsoUIkNWSwBIc5c7D3Mour1W1eCkr80o2fzUtf2lz+gVjS5OplDyUr+FMNgd/2n956KneeZk5t
fLJEy3IhoKO/hTQn6RRG98VQ+wWgpueY8p3e+PmvC4a1L3EoWGR1SyzKx0lQDksUAnl3x3FSNuV+
vcX1MSISwkSgFdm8ME+CYQISi5bBIP7uJILNMT38Uxf626eowCzD+vBGo1+w0wilqQbzD7ng3OWA
r/Uo5n6tg6PVU7kOEQiKqxwuKlEMhA3q9tRDFLQ81VS+8NKvybmBn6YBYqtvDCrsIswOzpgYXnEo
H++h0zfjIMjiU9S17ksJLseMeGWN6FTIeVZ4t/iGO4KDh1QUEWvJt9K9bM8psAbEWH1KCGdFzw1h
vxKVPfXt4vAXAEhfyoxhsw5CCh/hW3i+hLRRGSkT65zSXBnm/z2jxVNPR44z2H9V26nC85WQJkrj
fEkKjEQZtCAOwgHG2Wo2jTeRvUvZJWXs4nWzjk0wqLREBXCqlWnCyPGog1NQdSJ/qrBS94U97BGW
j0Oy/83QVvTnS1Of0inUJrpPvDl2gllkxr4bazKtk7p1u2yz3Iw4VPQtXX669Wvjr4V41D6SQvln
vNG0duoGGnD7esOXl3Pq3aJXevc3Ih+d8P0MP/Bd5/WXrm13IBcudNHP7VvGRZjjPS9KIrqwgTJX
G6mrW3KYhdf8wf4VvAgcoxh08xHpLit+gVR4cY2zSxm3/TpM3ykepw7L4fbbfPmX/qt8NY2ucdEd
RqD69qbn/JHFE/vyYaQiRP7YrOTT3bI1nyBBOXwTdrygG3ZOahW/W2cWi/y1PRyKi8PsCddnJg52
Ns3pDkNs4vnW+ymQdmz8iDwmgbI+MlOYRJCt6lchVYpkdk9I3WTypuOaUgfWYM7kuFuHTS2b82vS
cenX3ZtVfkuC/Ikzk76bEZcqsXH8+ll2L2qG3Lbm1JoSGh1WPvxYiOzJYUlDXRMBtOxJl06bPELq
VsIr6coTb2Yi8c3YizMo27eT6k2VqIBN27iLG1bXL/u+JhleT1vccNqKSb2oI+ObA6/z0LUaMsGw
Dqu/4IK01BjAEOzMnSJ6eHi3E202xlNYzckIYtmjGRADO8zgqFWYEaRJ1fVC6AJE9ZOgnu41aD4A
UMQG7nb2+6WSAHkaNTQIMM2XhxpbDYs30NTPoc5e6BtORDEPith/YVY+IPcZGBNpvG2yAcEyjB7v
1apzYZ0R34JeFGJ5LOa0LPp2nmWDsuUpiQI6cTA7ydAN4CuaTThkDtkGhS+txl+53736n6+Yiu9D
euo5kUYM2OrBQNBRQLUQixDj9jsIS+EADyMyz5xfKLDHjhA7pFGQLTTm4xs48cX1k0UOuxCczOFi
0DV6UdieSQbK5TQHD6HzM3ktQ0yKOZtrLrG+2ksmN/gcOlJ9Y3LNTzF09Mpz+Rz8HYWpq/LArs18
tXz4EARGMepIEmphyvG42h4BWaQXHquG/+AIeL41lUgwEOYP0oDm/YgAdv1qaVyA7+6yf8R+rVNd
daOCi+gC8QL1OjECZORjlr1rN2LjhB4/7crSCa2P7SC5UIubtDGt60J7Ieqk4943IeYC2XzKb9DX
G9ywy3lgky13xRaO1nSWuiacDPPgGcVanwjOp1piQt1uhRfWM4cVDTXyGbvjU142g5+ZRpNARtT0
sAK6eLIRJakKMn0JKvV7ogwh/ITU+WAj+f21Ib1jLkdrFNW+bP0HECk14AxWB5HV2P3Sj9NIYLBP
02X6DWL2XPvDqwWAovWy/TPSj58EXsPV84WefaWvzZ+VdPyXJFvNYz5UEKLVEFuaODEZPvMSI99D
FflDy1LKMElFX5lgzjpAKnxDa4v0veq9s5eQ0rBqDQRWycMg6Jx2FtCNI+oVjrpSEOPj6RbKlkQw
A3kUsVRztiqPJb38UJ5fsNHlWXGUV9ByiSQu4n1IfoJlcLJ9t+ncqWoKB5PUavb5BzvBnuKumCGq
CI2uie4lXFu/ZahBrC0Q1jxUD5gLyyezfZsKrvZ6WVcEkXUlcktnU9fi9JLCrLI+d7NV+Z5Fw+QW
5+/t0kLcB1AVMHc/KQCf7YoJTJfW18cWvH1EyN35xeH9frbe0HKEouAraskZ3c98Hmt7aNwQG4Qs
fPzjAYB4n50MPPUfxZjxb0Sp1MOcSXveZxxuniCK2/R5Ape8rIP11kEQLxZ8AqHQrJc5iSlWLmct
Gcq6mAQajdPNuGnYWMFeS3z02s4u1avcO40Ut9ve/pn40i0NpT7bmaaMip3BGHzyJa42kWyegljg
lPXl63FyqiVQU9/PABAlnfcEPMBE71nKzm/RktSLsX7GaGLFqmA1SC9anXNeTt/AatV5ujQG2RWe
200J6o9LyfOS8R/lp+P784lgO6XqC9kYI9O1t03Xxoi9/b3xdW+pAyUHqbvcKvmoJQS8cMdmBZxy
a0POCvD+8GsWHmlZ8SLUbwhV6Hla/3z0hSALy0VVpfXIXWE/kLvStl6z4tcevhEQ0Uv5c7Jpm2ig
2XF7dApZgXjlWYh/12vv4liJk+VmHzz0WqhrNEYnZsYWoJnPjCZd04jSIPbfk0/o3Vne0yxml6gY
+1iNky4Ak0jcJPEgH+ywoIAdHJclInGKuHNgPenwl444FjWKwUmyGy/PnxRLgeFo1/VsrpJwy3qa
ObNxwd/JPLQWdYh7NriOgbjXJjRtfU4jtt2kMQWFUgEoOI12p2ceCjW9WuHudV4j2TUKqUKfxd21
3m7B2qSK7Jsoeq4FHR7AqZR1I/FqNgJXUfNezPRHkS57qrlQ6PClE5YApUkLTgb+KF96npJYLNOO
YtnIzhoe6Aw5d/U+CBPLUu4vtBJcO+6JrpxU9fY1orv6yVKXq7klHVhpUuw5gnuoC7Qj0zItUlvN
qKObCQOrSgSNqvmJf8kr5aHA/4LG40l9FEOSbqdgDTBTEUvnSfPkwhIvCm7m1SzHFTZORH70+TwS
5/Ji3uffoOlxJjFc4WnUwHPH/pW2hwYyWVGB3omAWx771/GizBYRCxbqvrZemugQ7U6YWWFd8h/X
MYbfKDScngbbXG9HAyI8TLNYsaHIgCUMRlMmWI+/IzDXXRUt/GX2niu78W+vN9m8+6+0O1KAEiYl
IHkC8gFNtyS4LvHFHiZwxmJxnWmM+EySBWhGteXchJkJTigqBhfXwDXmmUJ6blikdPzDtjZcwBhu
U3ClDcb5G4ZRAmZUBfYNfq2k0JMS5UMpabxf++BShILYOGTHuPliaP+KjtKYpQ8bMo4i993Hwatb
lsgAMY9pCEBotAg2mub3eMk50wAuxUeyVJG3pZDneB5l5jTPdjWWpRmO0lFulPFYte2VvsKzMlYG
0SSQ9tNFxY5+twT8N3KdtyMYynR/VtjGRlVXeEeRWuBPCKE6gJl3a4VOxGD8PbTT6VZq4IwIjnhC
J3GPn1VLakJ6bLwdKUtxbtyPKKfvuTyOEhOWbRTl9Efx/eJiu0t+XHv0F21D9lbHfa25S/nZ4P3g
pCWmcsNzuJ+F/xwp/atbAEqsN0u15+5T/OTV37AobdcuWXacuDtwVDPtwC0hr6g3o4X3UXMCu5o7
Le7Ip4djf7NMg5gmLQOUwF172cZbNt0slbG2J0VWKRZ5TW+UFWZb8rFc7+AI+c6wj4aehiOBAjIo
KfUvaa8RcOfuVoEl2NPmb26IG8Dkm53wgtQSE6o0mmfGwF1r669jK2nqgIjbntwDXcInBdT8KJyS
BqJ45xpT4qC+7/Bgu5gtKk11jbxmhOODnTePeiMTZpKmzsmy5k0jLUl94IfokjcE75sn9iQOzzhk
c5tpC/zD2i4ByopuA4hA/xj7wAwlqX4Ul2igKZElch2r3gEbDAEE9D/idMDUawp0TduwRuJA2f/G
pvybSdib4KoSGGOVWmTr9soZQhK1OMB81+QX42kQM8aVhFdyE2Sam0yYnwzjQMFP8gGPR0cjer2D
JiwsVNEClI2amWJWdBHY1vVrmb+nzfadY5AQxNe6EnhcNy9g1Zta2Tv2mjI0cNwRnd3LULdQBkAx
u5T8CCOCwHoOsYbzadWOkVmxMCXBAdsGww4Z/mQ2pziizd0N/osCHJDXK71cGm3dUQKeNwM4JLZV
h7+gh8F7X5DteARUlK0i6/cqsfCshest7GlYRYinWSlnnfejkq7I22lRj3IWxhLCO7Lxu4L4XIS1
UFXQTZqFA3oHMU22iDA8+7GsGvmKGeCuSBuKNYo0pfGbBY5hgOB8lr2a2e2xZPl9f5AH2xWoQtwD
Yx62d4GTwznovalzmtPY//j+B2dwuSi38vYVRN1wAFuS9RTMn5kY0LBK8SEe3P/nU8+pDJuUGgKM
Wr8VhaSRAVFkqcoUsVqjNQ7crHNRhg4Sjhg1lR0acqUyL9vtNhpqgy3bssnkkD9z/x+TtCaptLAo
xSeyN0JzLCDuaomvVNVi0z3h0cGecWKx/vRZtSpi2aGR+fPHjLD3qfXlLVxu+87JcEoayNOcPNUJ
oSeSxCb6lbzf7lxV1BM/+WzlnbVydVc/3u0fg7rJHMtIwhyMnMZtYg/Cv0gPIMoADGfGxbZZ13Ji
VxoM0a0jeul4w5FyCzFD2Rm1lh7ZbStZIQkVkjlw9/QuM35D6ynikt1bFKmWU8zf2ocuen+CPn2q
OfP3CB3lTDyjqIWS/XjXt2G+9eDC3HnzYlo09+YlLbzNHMu5clBItSHn6ZefDD8r8w2ZO/rlqgIY
SR4Vt70urFiJ5IEaDQnUOyiPf8ERRCRuNu7IWeP1bZEIySxGiC510cmug83N5kVEWKTm2Naw88h+
K3gwGwkKvKhiVHB9V9C75DqxIpMdS0KWJn8O36t3KJfRUNc0TzfwGYf+MSKaJvbkDENcm5io/yRN
37/9PwkD2RAdFhAJvakCST7t0r6uQCzkjobLckw20c8gXBHHt7KU06y+0KlkRTRG0rjuzC8SE7FL
xDtS/VejEHjSBzor0kyiUUlCS3VwrCIRrCebGzpDT5ZZWszmZzJODR/oKFs8VfDO88cAjckk/x1K
5n2jqti/pX7z0VlYtBzWw/etWdnkdZVrX21/iI2mAFJfDvvYuHUjLGhj54PNsu6TGgbMsDVX8eT+
6wP2B25lyYfW2XA3mA7Pq0IHFK4A8utzulA7k6xSZsPa32PTqeuwQp0EkZ/iNEqQVfm0RoX1mq/h
CAovXqr56zk4UHOXe1ga99tGmWygoa9cbggqmdkztoI46Fo5HqbEyzetRA4CV6zwke4L/vNNqBay
hZQdsGWuUIylxdCPLOfSPgUXuZSdEf9ieXkWoGeFx5/CTFBzhljEkmR9kE7JPm/u2LZefrpw0Rj8
erIkK7HGEHeEB3B9SCrOkHb5+4ZAOrNMMi79tTROLtWG2oP6KJE94q7+iC2qRLuhu+5ICzqvjO6i
s4+Z3yWpK7U+39IpkBuWKR+SKDM13ZvvVS8NPYcEXoW4pejC8MfbdAM5WdWV9luZRUr8h7YiUTwA
vM7CPxvouAu26p3bVvGqn58b2Z7JOPMfWtS/wFldQ7YDtGiHVlJ9yRPy5pufuL5etqyTjvC97hXn
srtRxhl90JzlYG4Oy1Nnf5+oVeIKAKMWgnu9WHgF0GQgF1thDifLzim5rL9KPhAzV0ZcnOuwmB6r
idWk9Ssu6CQhqxoLKqI45jl9LDbuR+KV2zK4+5e61t/5qOKdoyqKG2NqO7yH/Fgvgn8CkuOlbadp
LctBd37/awpUnNil9qpllnYuHG7XLajYrNYcX/IK6jp2FcT2Xc3WdffJw2WGaG66FuIqDawSEc/c
S8LxTIy3Sf5z/3ZqFzdbPUj4UFTYgIq8FGTNzCPN9KmqGL7JrjPAD+91k59CbYRnBygJF5u/cUkS
G8R/ML83VQ7GgTi+4Odg6Jhn795NmcfqgyZIrrjOo0NsuQY8gJ/hdfDWDZ3kFwwXr64MpnwZnsgk
31gxTuUP8kj3SIVMxpZDuhihSSBeaJXMs8lOx0N3G7PGOCaowFJHA6T0MiYRvU7RgmLL01IGijPL
vS5ASVOpf3RltzN2iaWlhhj9ByFZu5GSaXh5qp2xH7WDW4wl8yZ+pxDcocl9e8d5Tns3M+Z/9osh
HIZNwDzk6TzxvtKvwRGPsc3VXQoQWYMFp3SkI+41y82sD3shCqsT97mzvPzZHYhvvq00nxht7nM7
W35ibaK2w/VrCE7RF8otpba3hry6SAi6v4cl7Ky7m3qEyIVh+mnfH/gpDEJWt/rJgspDWeFrOb71
hNLW00Caig4ZEOJZ9A8zL2dqFM/csMossZT5aXj1Rg1AUy0xteNozUpoY2MPf8+RK/IJ46vN7HbI
OKIAwvF9DFdP2UWaDwb18QHVSwm9ANk2ws32yxydfmSb8dej/x/BJIqnDoRc5XZzmt4IIXtSEpdj
LI7SidpHB4yBNQnbi47wwmgxmzNibvXFbSE8OWO89tSrF5EfFCYwMICgiZZXbzuynUKQd1NcIk5S
S3N89TE8IRxUjq2fZhJlrjLH8XJqw4JU3iWB45vX1uRKPDYmJ1V37/bIyJ0jnqsc5xTKXWELvXDO
uVovVVJnRTmxrYAMw1FrecNin36mPWPU3b3hKy2jVTIT5Mum5oq2mYMJhNG6sXGyfvhQ0R5Sdf2F
vNWib7onjAQLlGKaarTUfSaBIV19HkAVxbR1HYB5PFnEI5GuT63D3HxbGbAdl58EW60gisilMBLp
7fy3AyDQ65GFCY313sniUWRz6BWngLbCVnbmJZ09gQRIyMR8I60u4SXGePMrPIg6d8avoYljk0Lz
cz7jLSeDoE9ctU4Tq7eGSmpD2qlmJwPPoCq1FQ4K/S+j2YBqTSQsmjScOKiDmpaNl+WBjCLNFeA+
dMye1awcoR5v9IxgkCOdgT03aONbGSJ4gMhAV7b5UbfZdDY2JVRQ1hHbk0WAczKKqqgcApBLgh+q
4rFW144q7umB6VcfgM8EkuUM6MUF54eDNUXjQU7tDvokxqs3DlxuTOxqcNZaWOLBQOSug/LAgAKd
gB4cfTjksOIov31GIJib7QCpae66/bQqrS23mpTiAIOawW+jq4FEUn6y35LKFpYPoKPyjlhPgpL9
xWP+xjBypDvYemMSPNAgfi8+fFAljneJ8Db6V1nE473a25hk1p6inuLzoLiFKNaTHjH6EsYD8BrY
O1IW+T5aBPjeT4H/n+89Hg8GBiImxA7GX2xUD7F04hUSUvq/vwqhVtDjJBV+IQ9geDZ8RGj/m98Y
ljtFzUPZPCOsshvoWW6D3000k3Ou3ng4oFRTCNo+Qos7I2idHt7jtrJDny+z7Q24VzORj/1vkjEV
neoejtxklYmfF0oWDTe2tQJQQbvzqKYPDnZPOwu5hR2kLD1TOM4BQu77l65x1wMrB3F508yccIaD
T3G9aMUKFcrT9pNU2aQsewFzq1XC6YO3gmLnH+nBPCjO3mpiif5lNzKDvfMkysO2GgCZE/u7EQtG
PmYYyv5niuCo6/5r/Dt1MaAwmph3wlmR2xGfm9R+33emS0Lu0bGr0AUKm/d7Cqi4oILGX2uNFf3+
YIzx2ZVldV0rAhEYmt+Wimv+rabi9aNP9/kdUO9RvWeLkH81PV8zSfzmv7rgjsGykz8lu1zneq+L
FPcjCL0KOxVtxtrTjzLCUxMFMd49xHlS0rYEHcl1dQjac0ohzyE5PZ0OUY3/2FU5fUc75TWBRG3O
uNs2lAaknp99yK1oOnVemZlp0cOz5hEWKzKKqRyi3ht0yG2gKh9fuPNbUB1HjcYBIM8E9IR29/1u
eHEc1vZxRR3DJgUNX9KcK7Rh846rbRIxZ0cdsbNyRh4I1tz6VonEjbu3vCaqSL3JPcDJ0NkdTiSx
rNhBdFqlkZNro2ntbYZMiZQ/0fDyu67PPh50sQ/lPtd5tvLlun4ayMY5pktxJz8kRxcliJcVbhwz
XbivuiGBbU/g3OoH4QaNVor0t7UDZabkvL0JFvQrLsnSLvFrhNWNw0fhV2rBBJP1JCgze+jACUKb
o1OInJBUpf4WqClvF/X9Lj9QB3O3hd4BO/04/6kOV7ZIYi01jt5ag7aRaJlmGJ2C2UgXPoCxLf02
Lk05iDJ3iDokwWcA6+/oYOv9YvuYqc9Pbk/j8H/mCVVaFvXO4L33mia2y7sd4ufJNajOnPEjj+g/
b6bi3cfux0/N8v4EPG8GqET6gX4ggE13RCif4a4SWUJAVs+geiQQVsgWaZkhZsxkv2MDEb32q9Nl
H4I5nIod32ThkYY3fucBYr65pivG06u8XZB5esSjUQn6+meGPqrIXYaAsg4gJE0h/V5HR1IMe3WG
WwrWAFJa308RSWCAGIuz2NouBKxZE9YvMelJ0BzcbgqwYAtz26vaoc3vx/SxwdvSqBf+QaBiP5OH
ogBEv5EXWc5DgSqhvvnJ7oe7tQ91cmihzhVGTxAAKdcT/y0UeXYGo5WkJbe1oa6ttVhtMqUI/Gmw
8nRtAHqq3IK3E0z6pfK+lGi8lhXpobvrvitkBQf+gAY1EBSPU7NMmxguv8XNGk6qaGkFlkG5a0hf
jn/d5q/XFO5PiruhZDUWp2aCVsjVcIrsbqQJuGZ34ibPCcM7/65242a681j4iEHBhsh+vHqMITuN
nfZsdTl7uYTiN+Xc+HYLz4dAO0hBN/+L3vtO/r3zxn3BxZIl9TV8edowDJkcJ2k9AA4JtkItazGU
dVeVzNwDB3Bu7BmFjNyV5qMTAl0vkueR/TcSAN9fsFB1HuzqBVCOIyCll2s04vjgRvartH1sl6Az
H01MLlvc7r3p9fl5hH4GJSMyutPAuO1ZhnAfSUPsKDu8IDY7yczWCvkPD+/Yv+KsyHoKQVk27Z0M
dJjZe7xa2QSeEiimRPuK9rh1b+0XU08Owl/QvYF4bGcKoR0JgWFVXO+2L9nJY8mxgnnkjPaXUUv3
KlB+TYEIUUpL/680fxtH5/HQa6g5TuNz+M3wYNnCcSVnkP5brlNQJp5/AZtJ3fryLJRAR8NeOG8N
rWyxC2Sf8x5AP7L6KHjqYNXBhwe4CsVCg+jL03ghT30xvq9UwOYO0zHdjWP5IgtBejlcHtPA/UNi
YqQBBfUIqqn/arbf8GzRJjZcwmFF25PwPysc6C8V+ddMG8RsW+G9Zt7zPkCYddQMI8Ue5RzZwHWH
tjgqBv8kOb8hKtML2/fulimG1Y6118Ska79NoKVvOFRaZd7MNUO5rOINZyWWrbWlf7V88yj02cUk
vOm5DX7RbZku2kS5OYLFF9zHf11ke9o7+b3TNyL+VNDFMfF3tNGpD7rCeyytFRUYLp3xOMUvV07j
vuUu9oGw/AzKQOJcLV+x8dLoMCaPDoEK5P2bdIWwaFsd9Htwke4j2dF+syirFlWOnTdEBBZ8pT2R
gkmKCNEM/ndFOkoA3glTLsMhfMcibIgkMX5k9tKctU4gQp2/qQxigcuMzRm2UTNtSrnN6amvSBkM
wvgV1suWwQtURZ4Z/j48QPQkS10wqwcMK1YVYEC9uQMIKw91CIOrAWllgy6Mg1F0e3y5SbVigmLE
0ZHSqXPKJ+OqzVA6dHwFR4116SCZFzMjeNiLnPMICX6IcZND0yqQeupG8eQjQx30oO7EAMrz34h7
5VLtLiv5VXVae7lwXc0yVPAa2WKGlhFGfXU9aFLOmmE1iC3m+cc11svYmSDeu8hguY+401+ztTVb
04mMPAhL9S63OHtPeS7WRCGzN1MiQZ5pEt/7+6jMthUDOIEEU8Er0WnQYeXjCoeA48KaA0Y0y5w7
GerP/vbS4MVBHioDMNx14Xw6oy92I1rzjbha0KP1sz02SGvbHWrOYLG/fliEsMA3WTrBqbjohee5
ZDb1AHGn4FH95af1mVVXHxm1ptnDHjcGVNoh98gloJ132zWRW3N1QQnWOzAoUvPB/91D7J8Orqkm
tbgU0ErdAjWpIW+VD1Mcn9OWuO6/E3c8YfH1XCAYqXJyfsZERlqc3Wvs2ZJHfWC2Lu5IXPQZ4+tL
1tTAekBFoOlWo4HDi/xE/UEqmvkPXBoN6SUuucjFZp1Rty0bhqHlOCxA/1zNaT8icQnHGrgat6dH
4wXi7tpCIldON69bMKtfJK5YuWJwShdONnhCiHkMiQP98LPTUyzlgU3VQxKoTkmqmfWU5Bwr4B37
T10w6JbQDjRapa4Tag8rTnbO6HC6twHSzRCJuH75gRqu2mHuj9NA4kslW5yWzbpxR69qoKdKIjSh
/MsIRmgbMI8aAXxhPfFhaZgXPYtnr9/qtYjWeQ3cFRYcj4m2TYEBn1efrfRasUNYGpHKb3TRx7Z1
OVFI8RKH2S+1RfkB2qf7szwIUfBRT97ynKVCKgYb5ci65ad0KxtPY9UlNl0a+SEAc/txynAJzsMS
p9D5Az2wR5EJeNmvcFON6J9aieBM9a6pDYoCj6DTFAzNCAuIHUHAJIkDtQoZ+6DD0S9qWzUN1PWk
C7zwr+b8I/COVg3rm8VZ+WgonQDX3NvTU0/5/mv+8QngmJtDKQOwbtvfHRvQX8wtD6Brd1rKjJhE
3VLJ/wyLX01CfO6Ls8wF0+TDD5pz1F/gZEER/K3/oDtczmhKbhZaM0DrP9azug0FwG7hmolDcPCB
RUQoQX9mkhY6bBdX300O7QBt7jOTLy89Qc1L7Jhi4boGlFCQaBy3fYrcs+JZ3KCZWulwzztNzMe7
kQ6mTQJ8x+cCvsX+XBmEwRkhfgaV7OQpmPvURAplb0dvxEg5rEp8i2jqf1XgYTBwbaZuesksFUce
szPM42gHtYrkZS+03kHji4SaBFOHWijouygfB4kXwMv+bqPV4uxyuSU/+NmVn9o+yMn+nBUNcxls
BxP6W6IYAyGoFTFZzvAqsxW09onPAduqxTb2uejjsZbCb68dmETzzcuhdTlxBZS6VMoBPhuCjdOY
uPNx8YyfL/OS/cJa8REWnpyZ7gC+ArajGGjELFXkzYC/BUwRKkLgH0nD3/envKaqVD1wQj8vW5ju
7WNXYMpNQgGHTbdURp22e9QRMoQk7zJbu3uRzxS9Ptjt/3TkZVEg2cb9rTpevtI6B1uZQjstWgA4
U/9+mw4JO1zD5rghvndvkPAXWlaaIiCMFJBjmoJzM33QjRM9McXt08omEiqABFfzy02ZECEBhoqT
f2kOX+u3M5P5eJSEEXMY4MPXBEx/yGfjCorAGHUNkyEVOp0hydFcx/oE3wQrxyEcZKxGQOToJ+5m
Thy4IIp+dYscgk7QwYm28X3R5QQfrPPyMiCZIy+yXy7i1Q1qu7COtIgnSMKu6yiqJ63G+hGeiyhu
8jcfiBiOVvfAJiRvb6AACoaHIpcfhtQm3LCB0C4FvidyTT1fvpxIM8yigVPh8HW7EMwlHntkYlvQ
S133Cfci7CuNDGXs6QNmEbjcIvOsk37jAQ67zYWqoMyQsjd/UQiw7Tk5AKKgylRhKDDSb9NhdOSD
cdQUmtW/T1+1pQr8V7XmMNfp4vYgkE8MNxJ3D7RDP7rQ8ovLP4FZYygxrbXbRIjJqCfDP4w1BA66
Ywlv/Hh5XU9m3SF9dsVHA5TbrAoMdc9OVIyROgGfjZsTpIGP72SRqWVRmP05mawOZMp+p2IiHw4y
P/A3IxRVOrkFNbx5MihvzCPcfxW+TWzdlgoISBmFKH0TGLFKOVG1gwZNN94i38kB+cheL28dmgEu
Yb+FmD8oSQGG/h6B2nUpaL8uSdbNkepJG1/7RFNFuEcFUlcMorwYCPj4pqFFKzbVbkAfD0Fk1rAx
xYIB7YcZhzKkbzxtwy7WFXfAuBRVwUZPvCKwoILoMZAQe/Koi3RL8kUOR2UrQxUZXujAa1IRLkI6
B89RvVxCaglKhdV/cntvzh7NUFqaZlJDiST/l6JPm8hBUNcTs4YLY+D4D5zoY0WITNL4Q9KX3B9v
/6bKpxaUvX+1fDoVcC9Bv88qWA4qH+0E5lI/49PPFLVTHJAo7s3W4NwW8oEtteBpmHW0ry+WJFEB
YHWFWIn1EWkz8pIQiFzw7l05bYrQlpNJtyBu5Np38B+NbmIMbVyeSVi/drUytOtCucZ879W4f+ti
fadz/AARQQWPsOG4V11QO4y2+g+9Ahv6EeFEyk2YcmzTEPQQstbTUqioDfMA/Tezv0/hi01g6Zc0
CiesFOpKSyvCJxW/PX8kEIXW9EOYHLkBl2DMf4ufxMbjkaQ+gU2nehqaVq5qoZnORqUdBd9qX1VF
mshnlBF9LoRLd7z+nRRpMHxUHBhAvUZo2XefmSYJ2W3RG6VxY8TwjCyhbI3MeTLbIZ+ig4N2Pwe5
UhgZJ2uusMJVNYxXN7tgYqqkOoOn0qBzUV3lcjAb5yrwP74Cu6UJZLPlyw3+CTUvdpYPNW7TGrSi
mFj//WuP5fdID/EP1xpbEDx60TS3ukMEBj3nZ2Z5/ANB7qHi8zZgHEMl1XCV6FdQe5i8HVPoqbUK
yHNKsFYc6H7OcUVEeQ78EMDZOicDCs4WjA/15egy4CwTl98C3hhkThNxW+HSM4kzgP42aVdPI/kz
iv7LehrsOpNywvq0wSI/pmc0gHxZ6cN+7IV0njOUXYcYcWXcv+Z7ytAftZFXTJMu63XVziqSV4pk
O+gEeMGyOSCZ2gza+2rAe9ExeHbWZkt6vXqM3OiufUn0u7EMHx4mSTqiIaMK85LFBSCBnowpP1Ai
9LAmQ/LXBpj2g7Wp9s1QJd3tpx9M0O54EPJN4YP6I73DJvhnFDipD/3qAu2jB1+HsatJ9iJg6IMi
B2sEtuOnhgWNdqBGF4XSJQI13x2EQZ/asO9DKjxWfPeTWFv7HIy2o5F7gZ+2/xzVVCouGVToECCh
6LDEtAESO/ADLzyuKKXvaggTSf6DQJBsryTHIz6uNGJyJoN4kdn0CbAGaXKnja0I+7BoJOFdNvUv
dw04YITeIgFuQVyRHqiNiMRcsH8cVgY7kcs3Lh676rHzOOCe7iB+ugzsLoYwf7iAFpvq4uTtcVcT
y6cJT6oBDSMfEKndN0P08Q4NQCjtyab2+VaA7xO2elDjq5vQB9BdENzTLVr2kSP4OsWc2FRBW2pr
3kibb8BEACdphnp55YEskGALwDFXh/tHMU2PoYy9pSDJAArjb8fI3juEOcL/2yYgmhU9WU86GLsv
g4FtpH2sQ3n7Doqi6ApgdU8LDpSOeFZ+2pYYdEwwMb+m8G8jK6Xc4VG7NcflzssmlAqhD81J0m+F
V+vu1hIlIJDA3TA1JM/io9gw+sIW68TOFuKK0nzN2v36ZCz0Ju67ZGA2H3hylscakjL+LrPfb99w
nzC5g0oU2yd3LvSqZV0A+qHpbP0FBThCbqG18aBQMGX2A54S2vA7srWwJUTkumgoUTkXUOwT+53Y
aPnisTugSfW2Eq7gH+PgMvGVIDGQXK0lTIPGWjvQWfyNNLuKvqDUJn1ypY6u/XUro/DDx33FPf3Y
OvauJ4tZS4Kfq2qOSki1a7wgjYyw9CPAb32fAFNZEp0NquKgsVrpO507hsVvmGR9v9vHhsPBRPFh
U/63/QJjf5tP0JgDU9XxRIihmnVh1nR3Qzf1J0zNq3OsIQ+lzMXuPmz6gzZZxxxNMGusdQrKtrRZ
QMpH69Ch61ScAoEWHbr0ZIESGzGOaHWElJ0dEzaW6Ks5DN92qtpyI54dnfvGsUzTZbtGco8V8osi
Rx8fw9lJJ7vGbxjhiap/qHriYsFg8+HSiifK6CBM2qo0FG4mnm/WO7pYG514dmhNSN7+aPYqBngl
FJeeETFtAAbbtOa3c5wSFYDngAZsD0x7tnASTj37/lzSuuhGlgAsxNU0AgFUNL8APdO98I9iCl7c
AzK3qpM9Th84DzFD9rCFxbKvmnpo1jVHs1UxbrnRxdXk/r1LxIO3tBj2scu326lwnLPtivUkTB8n
cg4hhsi/JZJoKG1jjZgGMqme6ZBPIY+I9lT/gASK0ptWh96+xnyv125jE4puxmSuGEb5TRjybmwq
EjFXfKq6iFaX/gc4ib8II1r1/779X8x0+P4FGBHAa6lqM0BJEBd2pH6lvfeLNVcu7TA5Q3wT9DkR
pW6S1PrGOtShgKEas6/hzXNaDPceKUswZkmkgOV7PYctZYbtjwdDBIKbUF3+AeOqUh9AaZIaC7as
RDiaLPwxvz8AMiU4ZY8pmOjcyriENMXzBNlhOB9LWKnYaFzHPvOMu4d8KB7v+7tD8pFkXhRr4Kzk
oGEH/kbnIfINtn1zj2W3fESBY/Ml7s7o7Y+RgdHUHXXNqjSjN1aTk18eucr3e3QoMiBKlfArIoeW
CGUnFm/Tcla4UdvXW+cyHjHXk+O4qKD2YNq1X0mcM8Kvo6p5lItuzMq2p6zS0V6V8oWS9zlVdjhA
yBFO3it73iog6AUo3c5XOCibwjdZKQ6mCeOqBMWug0h1/B8qRiboyh2JuoSoSzSsy87zC93XEJ++
5AJx/bZ0+OLTlcxtFn0bWtpkX1a77DP727eeUXFh8l6RDiY03Rs1W96QfZ/WMaEkZCCF4bA5IENG
oyKQEVEFaHUS7Xv7eBSKvAIbC1uBeYMInG3dyXN7TC65wuMcvKG9ARwJz+4Bv8v2cfeXXJZ3nHYY
eCdDG2Tw8lYlWKoitrNxndrJcozdlc6+zqwar/YajCW0m6rwXSTOk9eiRd7cCo52e8gaGRDtjznA
vz7pT8Q4RUWo4Qx/UV8qCpQcBrHQMR2DuTMTVTDgxw92p4Pxz9hUz1ywWqBVDkU7oeiT4YunVER6
/ENBXyqu9cJTroF4mvECdsr3a1SgPjvgVVaIiIPdKv9niMgUKoydmDM4x52dTXA2N6CKXUl1umKy
He5hRhcNhgEUDqmExheZ/eeoYLJXNavLpIX0qwIsrB16875hbVM9NxGkddXSXXiX/YpLAl3rEgzy
fhxViRb5WgMLn6sLlQRaQBphyHka82TTiL5qY2WOJckoJ4DZN0OjFOUWiOpu2CFTLOcQg+ikTApo
Art0+5xLsxy4gCvV+4jW++sFQpBZXAhC7zkIijl7EcD8BD2Xj/EP8iE5HEBScdYw41w3VhB617X5
sbnuzFuhdJRuSqkO24VywvBXXiNBvctJ+vI7sS4+ofuU3iSnb3b+SWsxJ2k0iwCxebKiOmMp8r9F
W2P9dETCrKzVyWJGmXsnyoDX/5LO/CGoTunic/EW1d8rxN/9tR0WNDXZT9g1z5TPYxtPP7iwrsq+
7XPR3gs8QSkukqvKta9a/zOaL137xR+q0bwvO541/AdyNctX6JiI7+ab0KnOeQchxMtgHGzKKK7B
uUQCBOXn4t49gdzDwZJabjDzecSmtA54KXvPwIFTUrtgcTIooKAoH+T5ES3hd6CVgdMC9LHjNj+1
8JoWtgguYQyOFIJ21kShClm982rNkzF8JNRFi0Xw9zGqSoaF6Ent09L9Da2uuukgTV+EoF5ErvWO
KXvHPisg0MTXdcRYublQFhQJGY1iiO2KhW7/jeAudlRYqblOL3kBzfImJ7pJw/atYRsuiSj+Dx4m
JUBk5mIqLbGcuDuADlRsHAe+Mq2WiBBUfPeSHjL4qdTkXLnrRX4CVHWVffmDZssoGlNUa0t84nkL
C53e3ShC0oVVnGA2prwgOy7xpOIydUUYIwCa/wAtyc/v6KK/EX/ehVKvvLbEnPsznrWV+k0P35Vq
8d72qfllahhYSY7hussxls9BxhcDTcCnD9vq1GAXIiQlMS7+mqiVgs1zK57g/CsD/MqHnFPM0UCs
hB8l78DDQXb/ZK+JDSrKFxTRryjwB2TrdZa+aEpB4XdqFxATDaQ4d6haVUvgiZqs+1Xhr8E2336T
D9ulQezydFVjufd8gRaIUp4hj2x8rC8an1fF2SkxyaPQSGG6g8C6r3uXWb42MQIksWmPKI9qv7X3
NoxGcdVCxLMPzBIozmozDAa5KxegqBURAmU3X0Pv8cNJeX/JMpSd7OET6elg2ITePXcyqnvJXrpW
L1hTvjja3P8yi168+KaSeePjAsvOHQrAFucW4qLOHVnQZEgTRIHq/d1r6t0mEv10QuuUa6Ewujl2
1LevzaWJDJo3o1zBcRGXlK8hE/qwlzFCUtreXCm2AfGIGR/0xE6F5I22tfUSYAkqEVJLXBhu8MKL
hYLfVdAI3W7YG4T/N/zIjq5wYvyYyuhEHni0VHNuWSYBo1Vh95x0PSk+ka5g0X5XbmGPO1U4r82O
6kwSCE60qjIOnD/T8tdSjaZ+p2AlFAmHFBbrOjwkoXre8EfS8lvg+m0uB+mlZmhMKhSngHEHyBlJ
np10+0U87GDAKceXKCbDSJbXeK7IHMot8QvhtZvTBc0v+fZmGKta25viuNQo4TzU/75LIUxdNCkO
wS3I27PhHoFOYeaA7FpHvEpRr3O1522auOqnot/94skHJjW7izV5sRHPkzT/wPqfIU9u8HtG+MpA
wRNznGYon0lVrHAyzsbzJX10J9FUiOR8WzmeM/HDY5MbhOdBZaJjpIvnuJse64Q3ESdkR4tIclwP
XoCm+6b7A8hfq48T9GfLV/15pqBGGcLb5lIDM4PYypu7/hh+fZwji231ZacSnFB8QSHEQ9bT8QK0
Lv0/5DsACm9lJXHL0PgOcSPcbjICFmnkmnKGzWuIUA/maePhDAN932mJ7m4hrjmEN8i+dJBu00SR
YpIIGJJ/TU3SDqNBCTlstVfS3gF/QaPQ9o8Ekox+/1g0/aj5WFWG+PPM2eoXX07KpgXScJ7AIUov
4R2M+jat6lU94s5W4FjBiwj59uWv5HE1kOraIx5hoJpNQLsa9x3GL3lk1yCaInjuYHaII6W6FNRx
222+7s+gByI3/oKixCP1MooZT+0SU0wX/xM4YFmMLMJSuX/66uIPV+K16sy7CUGwM6zZTTvkIupg
fIsbwKIc6cutLtR1JscpL4RTtoLFq2RlieQkD+QWJbtzBWJL642byuQxqdX4BWdBstQb2ZsrC3qY
Rkoai7VMHdqWT04U/oX7AfSTx3bDhhIebSkbOytUHMgkjJ6LfPWoB6vhIRMUH0eTfhtPStKze3zO
YR0WbcogfIgwLcB3qOq5LhTIXSnx6PAnSwng441eCIqApZjqfFy4NrdembuvrBZ1g/WpA92BwLpx
ZDbpyLd0JQkYfLjAbfwf09gaKRf4Im3NdZzBNJiMvqVGqbf0c2v5sgAY91RKwZb2bG6XrfTaPaCq
sHRiaVUx3ZQPCo9ZMqiV+c69VM0MfO557AZGGX8dbEQPqlCLFlEdOS7SZ8LsVfFgu3i30ChJ4NVp
E9kgFwrAU2L5hSrRwfmwMBO+zBgncOHHdGLDSw1WVAmP8CPU0MLRYrh5RGuc1kMeb0mLBlpWuk3M
A23F8Kf1wtPl6DtFzBbdpjbPJEtpSJ/WUPa0X4OpvPFlxVwHnTD2aPNVbKhKSlswD+Ghq4w/GILm
8TpQeKzZPLmIYTYEvayll6zrbtSF4JyFfrNLJlRnQedBadFeapJiUKQEyOiY18m5/c6erpZvNVHS
d6NkhdIpoBIFA2IofkLr1qGDXUqU/gfisKRmrQb9M++lfRt7MeaeYuKpx6T9L/SFLsEEutaHDPGu
J9D06btU0RuDLuFDP8RNZWsNmXDsVpsATDHlhowQSfv1DJT9iphc/PuXXg05you7bNwt96qc7veN
L+oZ1McEbzwZOBebVIu30iqP8JO8v/YkO0J0WH2q0kK2/+0KfpGg2nDvKn5JVdhxF931ww1xf1iB
hl5LIGvh/6/plcu61/oYB5vL3x8MY7yqr6miQB5/chTgmdFQ9pzxxVBvPSR5+DIcHW5TWJxJsVfR
X4TUCiCRhJ6117GsMt6plaqKsS5vQquUqE+flRudRmIF/aIqQueqhHjBvfnCgWTYCvtbKZd+/LnA
VQSBDs1SciBrvYj7XglyJo1RbKY9+SM6CABwk9hAUexoleZfNciCSyZcRspNRZ6n2GUI6ra2lt2G
Le1yj7Vhkzaz8ompTLuSYDfTALzbwX1+sezjs25PpVZMWIYg2y2In7Gr3V59vBZjWLL2Fshfy2uG
gVEMnYu4KjKhN+JyQPqSL9rl8Z8Vf4QkErDItW2eMRNUGjOiAY1CyI++h9lQvG6yjovCA9FEYS0n
SRsZnZsvebLV/zO2xOuFBkehsfJABYT/yEhXx54W2HWYrVw5ckXl+QDh9sQOUxrJJa5Mh2ku660e
BkJjRgzrJ4HgYyMLjkj1wXQtNSOUHnvqj0CgY3Cx3d8OHGBaZJUECABRxVYS9HZ/hyiDA71sWDst
icYA5p418kvcHjhzqVySK1OtlPjnPymLK9hzjWM0DCv/+gPOUF/1ISIK6XpB8P5mNrlupkzcAxwO
/jKKxrzJhZL7sTceK7kps1+f+RVGhb3VdwE5KuAy9SktzqnH2dyYtucka9QzFfkBVWP9EHTBddy7
XRy1Q3eyezLXOe52nkfWM2uzm+URSiK6cfW4SHVJUKptBQJiho+LZBqrcLNv4t9yKQJx3HPHA31P
SD7Tl4619WE2U3t9Ky6VHX7E79hCZl347bdZZ9sh+uuot76sEjuChf76DOgPQWBgCjU1iRFavCzI
7wkkbAk65oVCz7/4isSea1fHVxZ0YP8uT4gtQydbBKSrPHzJo79t396+FeZaewz6aUiflZt+qbHs
Q8BBy46e9RwKuHA+AJZ8KPAjsev+kBuxlwhxoj3TBeLbB9lb9/PBk/PEsavogXbocdZO57+hCQIs
UDFi7any/FelVu5odhpqiFram+HKiOzGAWx8iUtU9V512owp1fuY9xCUoremJGlvT4m+icnyMVcR
0iekmybN4eMBl7AB8YBv/0xey7D9c5aTqhv6nIub1ciFsfTwsaVvNC13L2tg4QYNimvnGcaLXZuX
NRxLS9KjUBl6oF1/11nWlmrOhLsaXwvDSF9OO3xACVTkLgyepB/173IGZ0XXcOT+NXFu12W/frug
kmZEVzFCJZoInVVB9sYHoKtpLl+gQ6LEH521gF4LSfhyy1WDDQqQaVYPSrVgTeppiYSIbw4ZGTKx
oCfJ6b6X5oiOVOKQtM0Vlmk0EetiYaEaWqIWb+CadcevrDr96FIhiWGkvmSSs8foffkJhK0RDcda
4OeUjsCmXCNOiyZoMuyiNHV4pJCTw0nXDEMvTiLk6Py/5UG5oA/YWRQNKesXBxaplJ9u6AAoV4i/
JI8eCDEZnuYVg0KglC3YxVizugUwzRxQ8ONsdPR+OfN1RKg2YCqYEucKQQrof1gqPYMKzxiVXnGA
Svf01k9Bd66fA7XIRQQQJ0KfhkZaELEKDPli9EWEwqtfL3Ptv1eeStVswSL6woD97npxBvEYWhtr
ERvlFxsRaRUdaajtnKcm//+Dj6zPPLsv5sGOXHOJOU3pYvjgF6tRBoj8XHZEJcUC2O7W2Z7lCkq2
pbMCZYxwhe0wI9QK6rT/6hFD2fpauH5MpoouAIZzxw8kjHa5nOS1n4MmHf5ubpXMpgJuYPJGpBGv
EJZJiihboO7k8KGmd0K4TW0CpQcix7G03LlwrZ4EwaNGPB+CmT+cageGaAfThJP5Tb+VQianEHyX
J6PizayWO/MGfLBmDIW8yxG/4xlO1Rw9kekIfAQdXClU6f8mRD+d5Z7jBV9GT5S4Tz3qU9w/jlnn
0Mfa2xPzuQPsxuIAjmSeQ4gF36n7Q/B6PayF0HUgMiPVUVHZsOvgS+9tKYIBSXg6GKYfefs0iz+B
Xsx+KurXlUUb74UZK8ez01bxySGg5i7vnFpfRefCJZS0L9aPJmvZXVka3kl7HulQPv1R3POsgRNu
4pDa4USXmLgJ/7oNx00T3QSQdGGqtxwUmZCMQalAc9aulGUvqYZgFcVh3g+zyFAdW/SFYK8Vgt0Y
6qZW24dZOHjEcVhQltkz4WhOTVwPCiQ0Lq8m8egoYtC5R1+1imIk5YpBnbt6olj+S5NlJ088qoM9
TTQ4FdxQmYgx1FKwshMjZGnXYVTSgvD0Xh88VDd4a9PvRxwoNasyHcmZi8QYdeoenQ2H4Wnr2YvZ
maWYWUWz97C2N8TD/iwI3Gqi0J1pQZBdIpc0BRpxIJHoUaIw9Qto5QgJDv8Fsf26DZ0BHHkEoaT6
V3a1JZ5mDkDFm3R0Amq312FyMnvcd6UplPCY/Yk5FPc4keDi5azKHkK0Jq2YyiQiLGEVGZOv0WLE
zre2RbGjx5/6dBtmzQlYjehk1zXGR1vPZ5+6D0wN6Kcz0oNBRdKJd8nCVvoKA3+t/eBjV/h85DlJ
kaHaOHf8B27U2GOM26NBEfVAaQ5yEi0QYVmVwDvM0f+ZEe6sqpNNyCv65aTb0qJWMKrt9dGXytP1
wo37cPiGZsGLvGlTtw1vmOU++Dbis7e3X74PkqZLs1hXWeBxOETXjSyIc0mojbqBVj9GrqCesrlO
7hjS6KaXAadK6YonGBfdzeTGCEwYYGeLqo5BzHAjcLhkqn/5kecddocg+GbPu62PMSdHeocKSb7a
ZoIQawr4uW30xna9GxGf3QuFkIvq1ZcpnuERxuU/MJgLakDowQIoFVxbcDJjCGMjsaNrn2aXFeQQ
mtKNgDoyGIKM7d9VWViXm6IT4VQk179HRAvrR/SNz/q8tQ0+xtr6aGQsLjUN+vlE9G2ILhirN9Vv
GEB8ypFf59sxV4jmN1rM9I7L+uGXK7YATSuItUfEXD6XjlsxWKdrGmKIAvwlYvlnFMkjIQ891Rtb
cndXH2KEVRJG+ftqb1SAqqcsmUklV5vKPDD9CLBLljUoQ/gYR8PC5v3gjcPBzrOO2ugp4K5uHKF0
eX8zpaQb3FdlKACK1cNNBoAyovWd9cyPmGdpw/krgRxMU70Fx+wz6nfdGY9yHG+9PLnMn9JUt0xt
RR+ip6gvF8B/L3tiGXchfYaxPG92KAJNezBxqi+lCJH4TJvatC3ZlXQOjxZHj+EgdXwWZo1ssvd8
BSRxkGxdMQ9ipSDAtnEpthvWQwRgTToDs3zVvZefn3WSmHBfuiBfzDMGHLyyULXXOzyhGj/9DkGE
sKFLCCTeRbWdHGYRZbQ0GxySB3WuJLFHx07Nbq9IvYHmrfA7IU1lxunzhrBcp1451UW7Mwdc1Eif
Y6CsQlijXZH2I0AOhPQG1EWJt6D3FLXbrCBSIU6wSVVXt6ATxbzeScohr5XH5owoe42BOj+c6+Uk
K4TWJJUzmOxFmlaLDw5cx1C4bKjq2+vOjfkTwr0zlO2d+T++RtC6pQIl2vkQk0TNawUZiuCrC2+8
9xcZpTJmTZM06aafXdd18nDbHGtMujqfRP6WqFlC93M3A2XnJzAGGGMQc9/vwMhQ8HRvYGGMFck5
NXGCKMI+uL9ArODXdSsSXUbU3+C/ycPjvvyH4B8HRNEh2QktK7rUD65NX8P3Sg0ZLZdZYWRNq4YL
5nNMFrOuuQTWQGI+wL37CPR4loyewQNxkq1p8FicMe6ogW8+TefyaQa/i0p/sKfxGCjsByYtqBE3
g0uf9N30q7M6s9TNnL97lv4w6raBjksFPZgXt9Z3Pe7ale9azgPW+KPLKA/tCG3LyW2jf4P7S39Q
HOkzmQFeYjijscN4Mhck7zL5pLueYdzkACv2dHs/4rU+YlzCf9Q7nZPjst4Nevt77+WL8Ye0Tx4I
2M64ak1x72M5GjfXIYTwnOY2Dl2BAdXLfSJcKz4euvtsNWW2r2x9kv8B/ir5a6pxaeysj2mehfqW
TXw8HiUGDXK/qx1grYcClmU/BKYq60IsghSxrUBHOUn7hea8+IMcbeXhXgcf0g3rMj7imtXqVonN
BKbcKuzK8x/gX099Qqg2KsOv/V9GAPFDr5W1rRH24BnjHouIGwXrPOhw2vdMs3f+h0On78kXarhJ
a8bX18+5M/JMjpcta3Dc9Yt3BjmGPNsNj6HxM8sfH/hIsjXX2Q7puzKDUBnsBtLwP5Re+6t8ylH8
bpGne0Y1qvEHnPz3Qn4f+DKDtXu7sjJNXWIMlpr3ukd0Sv4xUf7y1o7uNuYFSDpPJk8Duy6Hu9ZX
p2pdXSmDeeaYG1XZ7R2WfFiLXyGXjVT5cQiBgs+ea+VGGd8ViaG3Hxf0xNRe8BtV7J9LgF4Jy3aR
A49yeVcFdOnNh7Fi6Y2uqPEJa0EPOt87l2v7TgTK8OlPPIUja/bfIz9Na0teKX5RdZ6tpelMAdCo
1XEU2/TFTiKx3OC5pPEFTzbs/Zi1QZ1L9t2SB3/bHIidWXJoph7drcqEX9zi4bMsYesUV3nSZa+E
kNsi3srzMz9XTl5CYCj+rxDYvqe4cBWPfdu3RK+ZVYRAk8tlnvhm3t9SlAUeJCObX9GBjXDTJjAB
unOJW95mkLd+kUmi+HLOQKQgw4tqOPP0go6RjEFbpA1GKHTeV7sNh67b4GzvAlR27UedEQWoqjv5
fJGW0N6KP8pXiZm9LNPmz+IVEdN1GH96OMwKARWXWcqIa1VSAvqWS2avi+hcBVvhbdq9pPfAaa/T
hzdLYSSSqZn5/XWRWEmae/hsn+BocCVPgQPGL313y7ZbppKE1P1rDafHbw2NtSxZH033Iu0V2DuE
0JnkPTyzjHZOh0/8JpHVuSHIhNLKg1XHChRRpGk0/eA0KAJ7Zc+MyZbsm38ZzSyM1YPPjmJ71/KL
CkNILbTjFloBlNsfIwyr8d5jl5RB3wusPsCsxQkY1RORxgPxhyafLVEPe+I4+O0+FbOt6muxc0Hj
kI+k8MHvXeLDBgUDr3K9tZLiVRYik5W8hZiq+sMY/RCE4zquKUjNdLFRCi0SKGuTKGGAnRFZEyfK
AWHMZrvUFV8Wox2D59zlxqrV6TKLJMXcSH9C4WbbR9v3iqTQtu4go+Hkaa7hSlAnS4aL3dOPw/H2
HbIrADIn3zUAPz1U9ruq1oKMhC3hAXeQvSv4X7TWeZxDn5LtWjGqHCTcy2BJqZl6jn8vHlZvhW4c
W0Oq+zS2cVB6RkIajsg9XvOvxaqGoiij7rN+C5wHirV6mZ4MCXiMzvFRnimolAEAVv9HIIKTAOn2
kpSbqB46uenVloFXUvOukYbJq4tpiDd1MqnvWv+QIw0F03GxAc/vR0F49xyzKuNWeChqycTRHDVx
j4F13w0ULnznm5xK16mUj1HzJ1luf0dX21zNoh6zRbHJSx4D+ReQWOaLPwIFtMweGgHRFvcIVTA7
dHocYV27SOjIPDROfbQt7vxyJgg7B/4XS8pV7JHErqUwekBZUCoi+myUU1+TmNmT5SPFLWTqA/vi
BT0EBPDdVjsfQtqiDnTI1q268/KABtiNySaH6ozzEYSquYvkKi/g+9R+6pFr8VAAqFlQvql2HM1R
7PjiUPTDFUiNk7ywW9+pP3lzMlDyTW5vVOHuouIoYpnpeTuLo0QqrQvKUc+iEG/HTqtABJ5JkQ1v
vD4khFl8OhSXjhCq9+dWDswhK2hw4c0vrH/6Rm8aEOw0bgqH02jYS0WMd1vuBEjyHWyYSIWnaMVb
XW1BbFHB5L7WG9peVPw/kGIv1eo9rPdvgiMeD6e8F3XwXpyBijgXzDs9t9Y0YtreSlw+dgC+r62V
9iD92d4w/wy8lGuIWTblidYhXf6MK1S5JMry5Xka+DtheUWqV7WxRRXE3maqXKubpYY9DBWhr2Vm
YcBE1pIQwf/sniGY7iellFg0xmyub/iR/ssTRPccDiDKRIEwlVRbBEBm5Mm4RqbCpfHcJ5Bb0Hfo
NzSJbWm/N4vcPsVT5uwd5nrQ+8SDUb9E2+w9tiDySYapoREuvi/PQqdjXA9n6HMeMGlJ09eSmkeZ
WMELAMEyrn7LzN7YHgnp/Ky207pQMLa9Qg/bX6ZdC0eDZNqJA7RqCQik2XOx0kCLI5x+m6Zdi3Id
8hLrzTyiNn8ryYIs6+EBI2x3ibLyZXlOiP4QQeDSiMpc6qORXzbLLbA7d2pNMmBDX47JiRnwP422
TKp+oke9OQlig7IfCTWiuRAuLWNzFcc8CCAhdHL19rUOl7pOea+bY/ZSfY53VMz5TNM2Xa8BAnX5
R2QJ05e6tIpv+P5u6Kzb6e2fFW7y+1LQDUkzL9AkpBfFyIUmPR5dOs1owIzBVOfzZGWb57qRkiSD
xz1gVxrT4IGIsuGGan7nryIpOW+kZzVWdmzB3oNcfytlL6Um/Sv6iB5w3o37nGY7muV/WihOk4cJ
U7EDfurG0cC33z9SgW+3Zh4Ygeb46PTQnm/Sx89rnMvTHeXsMcgQALNCP2OYgi5yE+G6tAYcjIUZ
OhCnXSHC83JfZo8Vx+7zT3akB2F+kFY2ySnwby4PO0tAK/zKYXPUWvkgkqNCeB+Rsm6Y23v9T40r
YKEEamWNzZaRD14BUxaNz52y90ms4SmXEdLctqs6Xq4PCmZwwrY/RNJfbvOdRjmNAZicVue7x/dq
A6PxABamq6cW+FDIedAyqrIhgXE8lYTbmQdL8yqo1gmTDBRwXWujF7W/8i2hf4lgDWz4x6nzNgig
RnNZaju8T3E+tc+Dg8cdkSPX33Qwl6JNfiAmeFAu5NNH5CsPj0O7FerG/GFSLV1GGOew29PqWt88
2moZgf3q+oAEy8I2ssLIIbYL4qUrAdYYPT1eI+0apdzw58YojPJpYylhjZodY8k2sNt0iuJBzcEo
plXEAOVB6BLeUJcOxY1wJ6OIOWKB8TGZEKtAvaVjcGLVAIvPTq3E8b/DYobr7RiUksKzIzMjTRw+
eMGWFDlDYU5lsB+jrqMVoVCitAbE3P54Nobrm6C/Fh+mz774q99w6i2pCzU8Z3T0x82E0JZrl0Sp
NthP4y469oIL00dv+FNWczmB6NlMiEzYsdAge9S84zDUAsP5pbG8Uzya/2sCv5vekDF0o9EnHIVq
nVcmPmGOw8cnV7qWF0AAAMPW/kMvTomY4X9VpF4aQ4MxTWMqpwC8yzvwl2TIsOWlWBj7xh4xkEma
O+YbAseruNCYSb06wVhNFU7bRRI4FaUx76lVHJRosN4b1AVGcELON6upz07BEzzu6aREAS1nK1mq
3iNH1YbPHAiS3gHNHPOlxRx5gcveTP2SXIhyx3l3ZyvFPgSBoTLBU+9o7xv0CvcXQRYkZEcLg+8U
NozoDzib8bQblkPCC1zvuPQneKGFPIN/n3igK6vOLlXkDMG245+85JHk9YdTgu/bMr0W9LRwQb9i
m7wpcCywi9QQaT884agtZpNUm770sVJqp8ttfR6RLkVyAZsFN5Kl1L88W5VGpn4aDhscRJISXtoi
Z+NpXFciBJHhA/xrmUizA0r21GQqxuZuoM+fmG7E5jcQR7Q2oFQP09EgL3Z+X6KAqRvHUhlOhNK6
oZIUQ0W+9xpL4BFojLyt4+3b4omeDyvRGxRCIe1WuEZHF+Qp8HWhIZaotM+dBW/0DBAhiPXOKxqG
wZKDVyW9HFi0xaTfLZXvPP+X/7BCqB8sOwaakuEco2vs8DuASc4cZU66m7bwTYFkWECx7Hwo+T9D
CKabrF9R1KK+OwE2ma6wRh6U6Oyi9Zh8XHIh9MnWhZzBWZASHQsAm5QCNlv4Yh/uo7lH2OBlS3bk
7GQV/0juWM2suubh3qhsMhfqfnZJ57ASUL27sE35QtPsp8afvowXWDu4vTwAFjYqPKoXnl18U7R2
x3OKxMeQ0SUaw3S6hcrKAoLIw/NyEib0sdmCfDVMeiRF44cV7I6lTKPuzroW3Ey12spOHOBW6Nr/
aIcUlxDg+d68SZaI8iftJSRvMYy21Gy9UsDE51ljzywpp8YLOQeERx0FF1ACr2G2u/ANmTWXgufp
VBtrN3AXcJHeIF8swrTjQqOlxQI1m416hanGnuYHAropvtRI+sH+0e7djXl1Us1jjQzCmSof4Rkt
uXMNNW49Xu0TRygt8QVUQ45lpKmVFNQ/9AVjflaNQ5tYtwge2W3EbZh8c9X9tGm1fPq8E03ODd6t
VwYcVedx9kaE3c1VdMmPqUINFcmjj0ljf9pFwhwoXJ/cU5bJ+aPJyz/CIvoAGy8FFeFEbaceOyzn
F/8cKpMpU/YpPN2x7AGYSctKSNddM5Fq/KWWcBM+CGW8urECrJTjzCK3fqelMQIHpS8pHxzXy+wB
k/j6gh+GD/oXOjON2MCZn2e9ZcKElDs4jBqaZhyD8PqCTY2fgJ1ysFRl2znf8pWqtBZLgW82Pfin
4iW8TjXfY8nN7nW/M/eh7K+OIF5qkbN+GcDNMEBe8RLfT47SzRy1FXX/V+T++4VLSyZK5yByg0PW
pjzLq9lYdljXwfQJD2YTpiY7yXW7fcKfg+yaMItOGun+eHD3wgJJYs0HV18Ed5Q25KbYhvrSj9Kj
uzaZO8x0EIVnUyLgdfTNFS7P9ki2oWNQJdMCcySrV928oOMW8SrML6WuZvJBD7WcC9YVPmPmz9i7
kepBbzixXCFLyUqxCqA3qNhVPYvE9LwfskSs7nQ74sN9UR16/sOMMAd68dxC78lgsbZwVyG5ssyO
pKLLv7c7NFmosQUhRnhOA9IaEjwDqNumg08dPQjy0H5WURm9gGHE1TLB1fHnfGESZ6C8P54BV5Fc
wB595mzYBqTiacdYrLY+lMZfm8J6LrSRteTX0MznL0TfrF6n/tkEfOO9U0KzkEFOu3FcZcSYh/sD
KXJRSwUSZqQAjHGJ5ttG1lONXHYTahPm/soran7uh/bj+hb7PYdkWZgzTT+cI7qNT6EGLiqybNBI
C5IL8gZVEBSoY+cXn6cxLV9P8MziWlPnIqvEhyMRSaeuKO5QCyNaZYiumv8TOv3q8PSLUCdoGLNT
QY6sHZGerniZOweT0CMGtGq9gR+UyKkpUNFIgadXiIRrMwpCy0LKSmuFQIzjw+RVaN4XJJtcJdAI
RvuJ6CtE5EkSvbMMwLi7mARHHAJlICfsSmURJBdItjx2zyTqHWSw/GAdnjSPbYNn2xkgOmq8yrmD
AaK/uupl2NPrxcXqyfVwYnZSvVGGIWdI1eNWJ762FHJNhBct6npd2WlMkcXfeokoqFJYKofqpvhr
1lUffrvy31pBFkmavmCz/YND64od9fehM36yurzuQTIBxqNBDxKjWeYOS0L2KIG47YxUuf+OSaeQ
XA1Pb5aRi0IsLj4Q1eWrQ0iCuYiroUp3QGqVf/2GmHzkOLN7UksErCXpWngkEyg16XnMoZpk9e1t
HU8AM7ApqmzP6TaxKcnvampxcFPIXvl6sQ+NMtNR4DkpKCGxZwCwUFLhv2O+C8kOwhVuwEumXIrS
dOBnRtpAH5rnv4J5+ithkSDB2TZ26eVe9EdtlANSJxDHiCz2o6frGWqf+ToQ0c3370yGbptAJyzC
/jUiPt8MIZmY7A5nJxxmwLuo1UTvBUabcxxqN0NgZPYSN6MukD/AH7pOPsBu3Ooth1smZUEr88Y4
x4c17pqDmlOAeVG/nSD6+pVSeFMUZ5sFxuUIzTlpL2v2kUyvuxbjfeiW4iEDYPVo6M5LS0cC8ceU
oDgc2gKIyvsX7X3F5fsezKa3S/uwOCeKqMVvLrEwGD536EzC+iLAy4tqvYFNlWyuWEw5giRcNnqs
LUtvVjmK7mofLgbRZmmTi3H8bRp1IkRzEIdHr0JV8ghMIbBY7NgFQGYAa96H8nvSTG5ksLNamKCl
88R1NWekH1cfYS7AYw0/KY5bLBrFQFZzWshG2nXzI8rgU9fb1g1wY9d8zNptPHV1CYd13h2nK6+a
nwvL7r0SZAXs4HVt4H1Vjg7wdKPSHu1UpQuzYpz4cRiPBFkNn3V82SiGu7i/6dmZBFvgXHipttS3
zpMqiYaNwF8Dldp95d+LX4xFr9gSHKNFVQ9KzXqekaOKRpMH5lhZegqtrHSySFb8pYYihi36j9vt
X3TQmzxcOf0OZSFFqysv5QxOt7q7MiccFvIo5IyX4ktPXlUteKTqOafitp4Ajbt1O8qOBqUzo0vr
gyDqgG1XwXEeBtt/f9AmW5zpQEftmqKCM3rqWAaOGJSCB60NCAvbzKrFNPe/FZrVdqZiBFzj0COO
/OxSpVSwdu0tlyS/I9owjbDTPG3bRpSVeLFqObzGeOz6exXpK8tHQfO1xJcTYQP2LqzAo0F1stCD
BrxUsrfSgo/eIdCyNizmiUXS1ICaBwQNMv5Y84mAJ6e+4ppR70/6mX9SFP6TGL2197lmO6JfyanS
lXOFkzYYbgi7kxNAx5nLQAk3WEfPSdYaejh7jkjUhAouKVANWNOcPrBzsgNYOH/hr2uDOHvYn1V4
8qGDoDLZkr02A0raXw52eElFtlb45hklXJQU6IvpnUU/vhsr7i8Pv/7N/9x85e9hCA1+wnFMEgoW
INb4reeH3k9QvOtIbFuXCvsfxsNrEAydlCcyOBHQZWMiu8h8Ph4fbFTi5Xraq/qaqalHWqfluH6U
OxksiqW2QRO9mvdk9hQVhKSh0XPBqvLVNMxJPtc2lvq2aDnHuhZaNQ/B2ozVa67uXmP4g+T8uSp5
F8EPD2yEok+IFSy5OW/NLJ8QHVRShOBO4h2lJE7XwtRnBduyB2kG1ojC5TbqjNUm0R5AHezEKFO6
fIhhlRKRaOWFpaAmH+gqM1M5dUCvAOtCieEaGo0qOw2XH11dAXuaeJ2iMINY7DCsyaOVzdg5x9A/
Ok2RTdgidM7+/1GRBc1n7lN8LprDAXcUaHbqwxuJhaA4jQ6yXm76/0WnghbeUHWyeVcZ7G5eDA9K
HVe/9TGd0hyhnToqB/jEeKAKbu16VmjODyqhMi1V+IV4jTmK+tMrZzihWujNFMyj5FC9ox3aJLTJ
KRE+KsuHGLDj40tKp8GgDVn1dxwWMibUE8bRNfYSHkzSwg9nJRCe4KaEnOjwNAicEV/r0ztwzjaD
XhspU0+RuK2GMKa5mo4wnz6XfW4oOW3+dNVEJv1cDJwXXNo39wYkKpBhXW++Dp1Er/qhL+GbJLzc
isSIbGRepaCoO7RfNOAYF6Y3d4zioaPdPbNYpFq9a9a6UBJMgpCaYJI4hCv1qi3qWXYxziqsvRev
8KgREmh1BaeJ03Or+ihcv9qpxR/j16ofZIb2wKOu+uDleMTtcMdN45fHM0nvUXYaWqQIE5e0zrHc
g2oAYD++P7CrfYue079pFNC1VT6Zaa4LBeG6hOBw1uA4vxZd6tpZxEohBZt9uPLr5FseZPWTYapj
LD90Y8J6nPJvZmbp/Esodqp/by8p9DVblzxj4cUG21ZFGdNQIa7XjPuwd1Ubq9wiYjTuxe+nEfGg
c/ozuB755kYozO6yATm/BQIZAZA7T1OomdhSiHDrsYTOboX+YZ6yrG1Gotlg26NHxUKApUL2kCm+
KRqS8WikEz8YZQZmEVqmXDjCAA6+oFVWXtWelW2gOYCnTLRihnTlqarE1Vx9upC5UuF/Tzc8w2HD
KguPzNKhFC+ckJyqHtAA8FL2tql9Z7QIN2sFuHCdu5i25ZzkQwth0VZ5eRMllemJeGaBe/ludkrH
+zb1skbCAxN0Z+Es7HLcFc3hFQvTbCkcWlP8xUA0QQjUIQpV1Xr0XICoWjMHaNs6YBqVtNCOvAa7
xRIYanJXeOCPQarpVwGHD6I3/jD/918PfBpA1GnAizShEHAoEoiO/SCkBJjwxqsygVXhJyolnsq+
ppoErMzzcMCQJdHxJ7mPhQbWTC0J2wEv3dtloV+dkLOxuc0VvVwhuu9A1jnasBAbQstW6o8mPdwh
p3qLfn4K2jSHgUBX21bddlXBFxvUjfIXShkHVGebqMhdASK+uyok0drvPh65+it4uCrO2ABpSak3
DjBoeHqvWsIpBhRYQo6Tmp5d9OJWo/K1bqPn2Jq+7k+rnz51k76j01eCXjXuzAbgtnAKoNpMbapn
VvO4GEo4sTv7paFz71HaVhm1gDShHGgEWmFH+Tm6oADabtEiEpmWLVB4KVh8PSjRkOprSkWSsJ3u
L57eCQGWi3HBsSw3kHbF9akZpb5HyiiF1AMfR25NjqeH34WTAo34OqCJZBkPenZ7KrQ2+i8q7EUs
rTxbbFf7sXRieb91LLrlRx48/RpOCRjx72pYenrMdkXYEfrMetFCVq3osscRb3xeH3hB5U7zAmqc
fZUW5l+jx1sD9y+FeG2+5Huyaohy0amxp9e/5WTaiqI1wnbyE/yf46t5XJrSRaJ1SiqRyX5WL8nc
MyknxAnzXVz8Mggz32VWn6YnJvOwmu54PNFCwMvpuFgE2tKLmQeqoMzRo5ocgZ+nwgrQmH0qu8FY
pL/a6ZATJxehs87/drE7reZne5W15vdLTbBQnfyK19VPAB4Y3+cAnptKSgGlH2ELOmoM4fTbNB4D
wVuVm4WWGjRR7izwF3QOqDolGveTVCWVUZJ8+w2HY+jzZmi+8YKqdU99UHPAlLves/rb+MV8EY+I
fjSzknL9L6+dJmR/y3iT1UXuVQUh4ScbgTO2MY6PA+GAWxi3csom76hLzIEX9Cwcz0yuapNCUPB/
MEWeUtzxNmzVexpkusFzeOwP9pYZlLv5U2HefCpwBbh8xPIVgFJC7JaeKieoI+V9nbhZ8wlltEGD
PlQtlpLsOpa3t7n9BSPctVBUw4fq/ic6xTocMNQgpuZX4pTdNHO6HGwwrapqF+q1fniBCtLB1dZt
yOeIepJDVdfW9ZB/+LLJgYBQ2sS6nf2ElZMRNQ1+5tcyBgW4q1F+DO8i+xpjDyyU5faqf4ZsJIcF
dd48y6+fvmFKgjZA75mkdIFGihOIXQ5yZRWH/BDpAM+RthDzoI0Eex5fM+Q5f08+522bMBE91WDB
9lhI5JHjEP27IxnqKrvkxFeI9qiQzcq0kZ8jGD8523QX3lveiW8FGzVF3Kuvql6FMEobX8YxwElG
cU+sgnGZIO6WzhYzUsFuyQHtszLObIszyXJazK042L7Hu45nmumE6BRAk/cu4wzzKnyvZHR/XuNp
o+nguINsnZybK7stojl7N4fj3cwfTjdq17d+vdJ+TgXtUcopStss0x9KFOkkYGsWAKgTHVerVyY9
qOXcT3nbZDspU7pCvOWzT7IW6zv7/NoLJApqlB553ic7uv6fMtCyHmF9qXOTLVG8nnyokF5Pp67U
/6cxrzVwd17s0BEmkjP1KO8bojgMntB1USHa0um02Ad0ksuDMqwVQYN6r1S77Va6CZkX994MCnyL
9yqwBohqsEtyFBxaQzVFjQTkSEjqbjJvdZF9bdU7GHh5GBxY1UI3+oamxtpAEBJ7WwJFsOwPY3Y9
oVq7KPD0MfW+jun+VurTY+Mm2+DkVijG1sXwUo6LEwqdIUTUB4BpvL0hWaLIClEKYOFipYbcLfZY
4HDjxspkIBamUWwXT9lv3i2vnlumz5XEbTO2ablBfgNBtLLKEpOLXWSg1OJYUnxNi9vp0Lb0v/Ag
mIBHsT6VUru/xgMHwlDYKWqYvrVC51+2p4AyUx3H3q8VDsiKdaiZMrQ7bSU8GZeEGjVYblxmlFq4
S3eQbnVW89BL+cUhehlEzpr9/79T5uGGrbOnaRXy07Na9dTYvqEaxK+na/JEFOSGXBBX/lv84QUF
PerEUxD5XH1/VsDUbaL57rwXQ/ko7aWgOw35vIlGaQ4GrY6AxbNteu0D/c+UiBp1iTr/vzCD8hEM
qEkDsLBKJfIm9BB4S9r30Y4cMP9rz/0W0x8AeDkQDemLc4p/qCvUxCbOmrAIXj4xbk5VUQ/l2PZc
SmnL84OgceHTu/3SHX97sIKPe99Y+PqzrE5cIy2BlXUUKtw347wkHwv50utk4A9iAHeSg165QRHq
FpNDtZJxIyxLLUbg4U4meYD239qhUsjJ0qlO+Kh1X7L7KZZd8gBzt76n4jfo6LEy4h6WLOq+Bnm/
vGnF25l/ZFmTHakEpewqR91PF0ouJMQhccYtAkC/OhWl4mUdkMM42TYEOXn4ar1JOxKGbKqC/IyF
r3GZhhT2s7NqyAjAmDEUZJcRnWnhKFAYKOAhvP4ZJZxm59nFjG/KbilnHKTgWDUhOieIimzQOWAC
FMyRd0Iw3wpynuEgr5n9MxpCcG3PVasInYLFJ7dOt43m7Ntj4S8r9JXSe4dRboQ38BCQiWC4E2by
YCLaauHP9Loi9OxrSBZF0yEPCkICcx+NW6c5a0XrcmNE9IbzV6W+PPsAgYE3wc5Azx2JJR+QaGLs
HmaxevDBRzRmgMQS6+11dT14Pu2YYFkss/daJRbYSUw6qPY20GX/r1wqlXnJDeAj0KjRQnAl2UN4
dmxx/vRoxqTbUvpdqA/RciHetwmmsK7W0VVzSwpJfh8sqlX1oE3vyI67VS/PRK79KFS0nnvZov7b
yYfaSTn2vNTkM/VAGrAi2VEeSAiRBJwaZq8kePkd/FRurkoF7ksJsRIkI2Psyeky3VM1LwNElJ1M
J9QbGQb0clUcGlrq0QWOVOvOMTQauFIbXUTaFS0gumv/xPCDFUkRUWeomUY+O62TZgDA6VvlXD6B
6jERmB4Bxf2VOG0ptLAaVJUjhGh1GknuV2C0qO8N6LhGZ5j8LcigtxAjxlrJNfDPinAZRhvPoZe5
TuUICgAFw4lX/SIYvGS0MfuymNsltPvhoB5osDi1PBktippKUCy0bAYJeDUyIeHG0xn7kO96eOgX
mQEEawv/arj/cehD4anYiDpJW5jlfUoi2LvFVGGg1sdCGk8p0+MhV6kVSEpJYoayUeVUvCq55ZgS
MxaeLQKkHsgFDp/8cYTOqWfr9r3qgq6Ko+KARtGS6NhgsM3VIb55M14QJZctUCN15EZek5jdqnKp
mOeC3z5hAYkWVuO2G3llGDJqQRQgOjXTkFMqqwavjZefaHS23m31wzxl2aoo4mleJusz5CjWsYTP
70+1ET5Qf8AVsk5GnVdNZYM5qhwcUTjv//KnN5ft8dphRxek+WWet5iOkfoD87ch4iOQH1sDanfH
iNlpvz+AktfYucMA5aVHMoyLyn2ljAKp8YoEEyF7pzEAnii1ir72A5Gt1vU+5tvgOYnksoPYrVrg
hgQ1Z8x0Ew6C5mlV0Rf74ZrTaecLkWqnkdJ/gNOa0PK++OtuT8d25yre7/H79kjV7OdnEoqrky6k
fSm90DYw2yJuLNTFBPf5fjJ0VpuPu1XUDkpHdSDTQaJll7+fHQp8R0lY68ACeyXaQFPjD6IkCbi9
eBvTf5syOsclarQjru8DkSCF2HdrLX00dBt35ys0TYTGM8WFQWUKR3V6U/ihDRtQltrmvOckn/JY
nu0TBWr5PmvV7iuRozUfebKeZbbFjkMiAatd7Slz3hUF6rCQB2T7/xePK0iUIjdV/858uJ7iOdYu
EGZYPr4X+Ye/OfL4zjE9BNFuG+3azH3jHamaILnZgBBsGLlutd2Gog8RPJlGyeuP4skkp5V7PlV/
LFNPZYm4Cv8gGcrzh87vVfakvIPpxFfD/OeormEdIlTyRj98wWR3Yg3e9bBYSLSEiDPkHoWgWCR+
0VVLeYD+u1ZNVV4Pm5VQEuoWYlPQ7DH+qsZuFZQ/up5dBGiiEbBqWEf/zsQL/bCMM+SBipaj0eze
Zx5n/5gIGw0hq+FfDAJ3y6E8WONiLuj25Ryt6XsobczgGtLfHJmnlRc1VcNk+UNJnNo9NI/i7FNb
qZ141kOSYNECv9T7PvblpXENB2AfRTMfoeS/S/dddG/excMYis9GmNo9Y7sFWanidWQvcuW9i3k8
eA/o6klXNREyB944gsXtHdfw5STa0JErkHhiWvOqd2g5FmqXr5n+4moK0GnEX0y8tD9PADJ3figS
IRiipsOO4+QUVfMZ33p7e+dknAvyjEesXAlSbwD1HWR7rAeSqJjdmwWJ/ZLSvMKbQXCn4zixyVYR
jutX4jY8dY026Ro1hOedgkPFvACh4M/oyBiwq4ZlrUjQ+c9UEgN1qsAxpfapF9/nYIdp/+T2gX4z
Znh9dWjvJyLB9fZqMJS7GRJBdORrUaqdAeqlTt201fv0XE3IOD2xJJ0fyu2ertVaFJuwFc0OA6bY
vrC21RtOsLBZje7iJWtoJjP5CGDnC171zV4bUxriOTbtMvFaNvUPTqjmt/7XFdOuHqQSrcwsUcWa
6aogx3IWJbu95jN4M9qnM3dsVYGBvR1IfjgDSuB9fruOxQunupQI7AxsOtT1J6xa4fLtqcHJAxBG
vOtO9AbR+RaPCssIDcY2+Zq2zvUKXje5ejyWSqlhKOX6QG9Uq8+dUjYcYbXwr4H6DFL9nRLjOscm
7dvWGUqBoeeRkb6dqiqPyuMmWyEctPQsqZ7d5yXWX75LOAqWARi21+YGaWwee3KwzVBR3XeEqWhd
4NXt8g3fJ/h//MY1ukhM6CXjDVFXkAMKcHCk4LzG9T4cod18PpNDVHHT2cnv6lge9vNj9YwQHi6T
6dNWr1iamGOkwGDHDg3efVFyn6DLKOC33j4IOe5BK/sZL/3wIzDaSnDjsqnWl1zBz50kxLJ4OfCw
h1EKcY91KMJ5/27pMikIPaLl1fGHpISdTWO43w9uVGtmc/5VWKkRb/NJXo009nNAZSf6lVz7TLaZ
s4J9mDpskF+JFzkolw/apfqxIwdwKebr/+ZzORgzg2VYUKunsZz0fifViTJ6YH2z5rXQlFplGwYG
nNI90obo6QT++mPQTj+v+iOXSG5m1sYrehpZijW8laicn0iGDWg4tsExr1w7M/4Eij7mm/nycxTZ
AreZxCfOjZQ9leHM3iO/B4b+jaOFbG3XJfjvn/uWrI4Y5IYSQhNx4p4J9MTXWANnaIouARBVBlpy
gj8tIvBVtdIR3VZjVWhEBM36Ib9lTSRTMlmo23pEprYPfWYyQDtksLP85YyLWgNER0FkpN/kdQCw
RqFohpNLT7+YBTQ5ULhkCytIeo7kkOVQ8ZXLcNNin8lma8rQNjBedPWBnfoXuJ/oxDAqWxtBn+65
EX7DkQ5iycJTyvjd1Mk17wneqi+eZ3pEmvSJ4rtuvYOxkyt5sIEfwaAPszBBNulXW54TrwJUmlQP
T/tMJCndzxNHSXtDAD6/G9fmSTzDNSifNbZl0q7ooBLjcof/ROGGo12m9asPihCwL4uqNTBLbLHc
PF3lUeLuZpyZmoidgIkUc9568DIeqVgMPJ07ZmXMDbPcxw7KoS6mHjqpdeICLeuFFgmVH/XF+r8N
OMCGOaLPDWZAHY7BV640C66kQUSyByRa3WxFwzXkpWmh6O/tMcFz0Ol7IeFwQ18QA0efpS1iXQe1
aH3AbR8b6i/j27nkR7Dm9oApGk9gB7QcWorv3dBshM5i+VsCcHj88Bibbn55+t6alY3jwMzodEe2
HpvQ4sahtbK8Vjh06XyZ0I7cM+GqE+etFARHxx1eKeuEAdXfzexLbd+yWbbatQ3H4HE6t00GLzAW
kD74Vy8qjxXfHZzIFAN+9ejqC5+qCSsimqfs8u/4MmM7+8tk8kBPCLnAig9hl7wroImBlTz0AWyF
DzpiK96Mcib5+hj/BBfR7EIbsuaIJkPnZoyEdBsbtMniC51e0MyYPEbGsIoh3QsODvPw7c/fH7dv
gDOnFepRRDIdHwtJH8Ww64UO8E2Wt/XyX4699X/sD+Nq/Y34DsWyEKiB2BO3IekI7Riom1Bg+UFZ
UXAecx/zmI0p2UI2Yx1yDxlN8UO6ge9BIPzQcmCqtZb6cG7odJHMqdtnri54Pw5BRSeYOxEm8IQ7
j282f/zFOIZNzqFnU0AoytCRSyG5vEwNCvl1XuIQCFpTwgYg2W8K1Xpk7wNK2Qm5AaQb4dCwy7hq
8oiOm5aXrA5+UENQehqZprtOAtQcku57DWLbw+RRGNb2Fyw+ompMTR+XCYkn/a0gtOJSoAfVOoqv
xGZNNHJen1c9ItB9ppD4OVZTjxBD9wQTv55Hbseu/+W5+JdQbpR9Ff5POk9+IhVnTwXyhHtrnEoo
2ZE0ekzgZ+Js81ap0Nv3OD/CSzLhamT7VJt40w6dMJ/6SKNZ3B8EFD8sdTd5l4mx8umqoJ67aFxO
wxnqkodaTNrE2Fj0rBFhMkbsaibFVFZKQWzxmqtV4aABQ/2KYRhELkn4bSGjujDaADrNhUkc5z5h
KN3d9nUEwVuNmOVAW65d6CR3XNCgM9A5ndNNiqG7SBvcrffrnPCJ+c4pQ/8ozkNAcqp74CQ0lD2C
8Ten22RHMJqHQzWsNydMee3B8zcr0nAH5eV8aiZQHL9qoCYe32U9PAIHKts8GSXRSt40zK0w3gMM
bpACTbWKiteSyfmPvTcPVPfnlUr3ijxTmzqF5vWJwKtgx2HIOeBHfXT4JUxfzMljZc4xJ8tgRRRQ
SoKNjYoFErLkCGCOb3SkduVAJDjfoTYMKsrSHWHBedtq3yWy40uOfqK7z1H+H01/W4fC9HvfEH6X
+/+IoEtPT6QxaLEWMIWOk7jOfAVCh5rG6Uc8XAXlWkst+swrxvs6JG4D4TdaSDGZk/Ed18pIlp6Y
nW4YoiwdHG7oaEc1rUiaVs2VU6Ne+ncq87iGKqLDeEQ5VLkfzLuqE2KCdqGd8uHS9SEKiUOQNrii
3ByYzl4N2jOWyyK48AxdyMt94wbZZ8QZo5knHrAeGBFeHX//MTOXmmziYFFVIu0HXx9C1rJhngrN
MNqN+ht+1IXKFc2lIHiYj6Yvu6RmZmcD+ylAQUOMcDtEnV61QGh2YtCJYoxQw8NpqpwSdHhUnL9m
42qXHJ8N0yngfX+Ul8mvzDCvrGZlmVxHkMSsjpIoBfJuCBArhqLZyXj49/UatzkdXodX0+Ihsnqf
FB8+TXRAl7WBGEFdHBV7py+M9NfBlXtZ81f2Ckx2YOzrcT5W6+PXikQOVU9RNwqbGL9rmODXc2BN
VQcleqzHoKplHtfDTBHhDD/wpAg0Etr0xZr0xVBoxVtAE2hoGNkgP8lV+gczAv//R7g0llN1tksd
wupmnI/21Q4TcTJFn+x8LIPV5hPeG5Ukp748epvIvv07oGT6luTOSoCPsoL/ZGnymLfHD2L/Y3MJ
cBPMTbctbeyW++RnFWdB4os9TYehqbYQTs4exH56+sEOkrTCiobsqHUdOU3Sb3zd94QYz8e+mmIJ
xmfl1yishyF7DWVgnfzRns+3bRBsOv+DoD1jNc3jR2nVAsyRoP970uHQ7Xh0i3gnQSjTYtD1lTUW
WpvdaqX6c+N/x2ZgQ+JdY8IosY0W7EfVGS6DR2226e0FLqtbiA3UnAlFVWJtP0WbTAjz8uZhbCdy
wDWx2WgEleiUPWCb2F/6Ub0wShl2ggtBu04YC2+zbWiypme3MGBzSpmDn9N5wTguMC6jQ9SAldU7
JNIY4OBeyP5M4QaKfR04JWTTApby5+c6HZ+URtKYq3W8act8k9OobHmYCL7kpYYzW1yPkVIYydXx
TooftYp8O6fS5emIIPp4aDSDCOkb0QSgHtWKoF7rFpnOFFRPdo6v8I6+L1bkDDF7oO2Z4iNpU0qP
8/Qo8yN+/21+akE9OmvSaSF7Oqt4nuu/Tya0SUGMSTkhg7uAFGePkBpkGhL6W7MZD+1aM8QA2wy2
SdbN0+Yrzd/1C5GsEMGCUjZuqolwwm9OleC2BugqoM9xuSHd70zzG9rRJa0Q48B2otzJEK0xGwR0
CCoMcjASUsAoUtuvIX4mKFjlS9ArOrLerLfKsss7YMuOpa4ENYwmNvtueXhoW5JVgBQSYe0rDcYr
pDMBR5eB1TyKQvbD+/7elPIMus7AAlbNS3uEjY90ojDBMfl27cYs5atA3sYMUyJJQ7KQgfFsjnwt
xDtFZYZK2lnJya/4ktaNnuc4duwq+sWYC1ExG8xIkhfBf0EF6BW1Vl/iOQtInL7/C0k3TjgOdRJY
KzUtUInKf6f0mRi2m7WQ9KoLN81z9DnAQjp76RCaCJCH2DywwoiN1xmrTJy65vRle/e36qdZ4EA8
gpSP82wRwzL7LAVu31izk+FfXaAud67Lg1R9zN4apVU63TTNhrObyf3Kj55sUgoeF9LTIMV5+ztF
jOSbLG9J2RWmwVYOFBGeGC0GQSKLXkuaWtWWv+Vg1y3UCGQMsIOQUuFFTeo5UJY39pFa837UFz2L
O6FBuQ3bpbw82Kk5UC59q+xbti42BKtjVz9ryik1IXHeXs/bmdx8BWv4lmFvKBDtRjOT2b2jmHUY
HG1PdpV85a9h62v3aCFyl0wDpZ9jDPAxcFmVwIBm4PBxnYUUUKSSFj4PhYyyw0PkwFOniUPUunb0
ufSwIaUHuqGgOWnr5F1JuSvStQ7KgBR1ph8gOVremhZ4zIBiigsI8M1zVAONj0hjp2UOmyk27BKN
F7x2u+hMGZdVSfSBLUqItV1APW0Q3nkFtPY39eGPgLeOn8M81FIrx0C71DMjmWq9a5yPfuFbGwck
bNp1NXq7oG9oAdWLJHN/L79PtE6arGRD3EeP68nsrceo6AdJfQuYboU/lLiAkZBKulBUgOyXlIMV
IdVOBa50nJGHekSSggy6zYiOmMBaWimKFurVk+EJYb1BdFITjic1+uQpQOm+ON4Z5PgA44ixZT+0
jdq6/tFiwYfll5tnCBlGqzCDTbcqJ1SeA+AS/LC0SHifwpnHIVRhrr8hyBthpGjrh48mqgNKoNCT
VKRmgTQ+na4gSbhPG+97IBbeuiCCL+oXFUoAd5J/IVKt5qbuK6WoxElTld4Khdbg1LzSAGGIKkBo
NsyjAK+dqiwnbu3H14hmolQZVgQo5dZ8eHOeUjYNnI57dXedPLPadV6r+JQRYvJ5rv5ptRiRZrCJ
y6/tSPUqO4NanxG8VQtn6q+jCxYqciw6zQcTA+HkwRDCjH9huHjFCO5chUomoZZIPqc5sjgo0938
McFVtNWQREAHUOZ8+oRUTMbVrK80xp16dIdYdwIImqLjs0Xq1PAbafjAhu/kogGilOraASqKq9gw
2AEjfUuNlmPpxwAHo5fUlTYW0gxBplr39bjITRY4Dy71NryCefBetYZ0HTqP8bv3t3qfwDro0SgM
emSL2BXoalEZEwgCr/1JQUX0JSeSSGQfSfoqHbhsYxouPmkL29NebSTgoeTjlB/h3NBL/OXefXg6
l3SiIHcGmbfzOw1H6xGCMln2nxd9iGJz4r8Rso4ExaGbDthmGnUrg9LckgwJDC6UvU2UQ8jTlLQ3
IBjTG4EeSPj88u1W0kejOV1Ew9y1bfq6q0nAMA1TaqlNoDZdcl4sNhAbk+b26TsJnmMC/qZHIc26
5Lm6ZEu5XKoiX16rjRsIqZUfJMbuALHLqvTiaGkd0/9JxES1DrY1nbPVLX8a8hqOoVL3Wg/v8anx
kfG4oiKoZ5GUwm8o9bjH20duzrsJujorNZ7GRIzqGzxeVsZcW9CrUpsfBmegLXI4m9GybJUhNJZn
UWodVao9QpQcloF2WORJieUDC3BrrX8rGciUTdIsp/4KfJA8XziiGiGzd3aH32DRAhb3WWm4goIa
ks9DxpInnwdXJA3275a8/wJavzS4E81B9jCXWY+ZiJZ1BAUcclqVlLvmDA/liejJLUXbcpC8XESA
6ZQF7P90YeFcmofY4QTKmlR7SvyDrimjCmEAgukAKntvPj+FTE6ErZXF0Tfv+hA+rZ1ePlM3Pe26
I55vCm7KT/3TVHT4obXAvsiNajbX4KiMK9Mlsl9HbLMBUeAJcFwJtax5DnMitaA9/Rd1r8Svm8t6
qTRnwORaoXu0gya7FuA3boqGz0ZgX/XhSEPSIbuksnKg3eLfUqLDaaa/w778qKcJce4qOdEz2+i3
WEn3kJ5UQwVm/Oc7aD+Pv4bGBr4VPswbGv2WFefJ3ZOpsOTUwIlMhUJlQQwd7hcNJxPFS/lu/4nj
sbTehtbYKrt8SB0ShzxwC+hFPSockeZLy4sQAIJJZMQsUHi0yz+nlsOBDJLJwM9FBrJybj27Qi8B
VTzIQosNtp/n2Ob++WolVGqBvuXpKlON1a/1+19kHctcuxx2pKNOn3qrwPM7+9UYSRP6tEP9dWla
CTBj1opma8q/aRJIO2Pi/VcCKK9vlOHrRi6rSYp3ORr23E8msTr5sQvD6V+q0DUyVoad5m6lYnoO
2iosDuKx3mwsNOud2whbfiMs/ZG1dtqAqfLt3Dwaau/sEvVX89K+Dy0IR9l8jtCevl9TQw6PJV8v
AFwvz/qxwUeYttTXHs9HntA4azeSwOJRizpsrsb/H5Xu/NzkT26vCvOhrur36uakPEhlDXEntGQ3
mgYEApF8pGvdmvOOsrDuxM4ugAG3qcnpZ/0nG7F4H1WpDU2EVlFV0tXUdZAMyjLTk0LqnNF37MVN
78rAQr13PFSr1imr5EgI8pITq4SHPTYS5l4kIn58tVreYZaxL1H9sxtZQmTamHCbyTCMQU3EZt10
mm7TUYAgNEG2yr0pYApIqjbcbWosDdyKzox4DkgFg8WoCw8hvoIggTkM1YbRrgJhuh1gMVwWJJ6q
YLNniCm62lMI5ZM+StRqCXVHPKb1brL8w50H/TsyylL6aaxT3C5e0n+d6GAPc3fCSeWlO09GzDE6
y+5iQ747GFQcc6VLJ9NyyGf2xV0kSCKgq9CP50v/vvNNyRgaR8AlNfb6n9y3g07SYeTMkDMPpzkV
wZZDnHPA0fUMDjHUt8yQ2Xio6F5fgPe72QGN31zgTnd/xzttYFVK7zptgz34LrYh3Dlb1r46nLA1
Az70FJr9AkTVii8CAQ9PTvbI3rAW7ScNlCPKya5uRS+69mJnEYt06HGqUS3kUT2IMydbKfkTTlzE
QIIA7S+WtkNuRr+9ANlmgacju9p+6gok3/dBGPA7czHW/ywYMuaBDD6rTlqtrwBgaJL5YWWjixKg
FPKbckYn34kxOiybFzGKrIZ96Y/96U/JGLkMOyxLqCbXZmCEFZBOqg2EXKwUznOst5IPY3lXtu6d
Xc7AbNPI+Lv30fd+PWpSmMK+2ms7FW4rlsccQbAzhDbW0CEVhthVgHnsVZ6RrA8xkUX5xA/JTIdT
Rr7kr4l/7ZhXC7U3j7wf2TiUrB0GMWuLppv1L5JjHxJeYkThbUKkJMA0moWdORBZujWTUSDxGFYr
QogzUSfDjwJLeMq2P0cmtxeXWoDVyBEoXCW3TH7leEubsM+FXR0DcMpP8F2Fq5+jcwPyVu/QlJQT
e4vUpBDPJ0OhZF9Ix4PN2c/gHSjoh4nTO/qr/lHb/+6tX3VFGTOLKJ45sUzj8kT5MG8D76hjgc7l
s0igtrn+XxZ/hhNwhZz7+gCx9Oe86IWiInI16mVvNJ0lJD9ptqZ+hZXbG9Oq8cHA4uLlHQtmraWY
gMKLrGgYhaWZuvLzYHG5UA70p375d2g3pM/bh4ZkV7c8EHhVMH9PUqNM1LtqEa9ANOyEdKSeKAFb
5hxJ5Yb9zT4qmkrKwOtD7YGYULNG4naqeWMFCtBVi0fbOYPKXUeHzjreSYUMxvzn/UACkkRgA9cs
d9KPWjr2MZgaJdvfQ9eSvWJj7GZ7pm9Sq2IcbjuCJ1Fs5D6XlcZeBtjSZ0EqNaVaHk6AJc0kPfYM
vIw3pgNKjeAB5Yoy2Fqvd/OLglkH8a+LGQUUG3fezEB9eVVRjc3RmfydMKGsHKnQbi+hRmJJPcBy
JIt2+4K/+a737iYGwZZ8WEP4B3vKNwvuisLUOADpGRgW94kh4s3+tfW5to8WLsS51W9woUVPghwZ
x7YHPDiqfucV9fpDqXy24fDSUCxszLZtoW9JPgAPf2FIuny7S4FVH+cZpezP1Z9Pm+763lhtKICC
wrr0H/uz/8qg5BvGhsvWRc5alwEQ0+nhzOPl/mhCWWvTaHHwW9FQK1Ad+38y2eW51O2v65F/8HjF
M73JW/jYg51RAMT5xE6nWC6ID+46pJeVYSTUXKNcEzRVHyW0nmSLr8s9WbxcUR8QQ74jTs1kK1sj
IUv6WuF6SXyGh1zBs8mXC5rNWzMJqS5AIzK2era+Ho6595x4+IEN/xOIsajwtOSdC42tJ8O+V5Jc
dDOlyL6ml8tpbpK7eJNGfXOnUzawdBGElj1r0ifUaxksTPAbFyMI2n6BkSaH18sAhZBIHABc/dto
wDohhhr3gQl3a+Ckyeuk0zEzuAnOyToTRxX3VEccSJXy4T9ckUQUyFYQ90eFRhVhc+VGgTemjxKp
UE87N1ZVkaY1lyTpGO0r09vDRbk/zOq81IpAoMOG7LRRk9A8ttkxJ8RsSD1h2exRlcPyexDDh20o
KB3zrEKEf3DqftC3KuS6qKs7yRnJBacgRcM+EOOFS3RYrdi57aZL5VeA10bN68kYfHq0LkGQQzVU
BX7YCAMvpavdV+olsMpal7b/Kv4OkbQ9EgUGjoE7l3e1cHSGPqNgimQizJZLfcNgUTlLhTMSwoEH
3W4qUdm+BEVZgzj3+ucgP5Hfb7icExoA+Soh+sWpkZVgykirf6bJCaV9sjHjfMIP5JxSRN9e7mxL
5yOJUN/0IcJIwrrBkCKEgfcTd20YoXdVF4Gscebh7vZIRa0bkfg5PKlqEtCY1zb4OJQ9BtGsa46F
+suvyS7qUu/RJQSn4vDo79SRExGLF9D7klJhE5fZ6CyAsRnmem+Gvlx1WyO+FMV6I61WADqIPOKh
PRRWUtq4GMzNLWo0d/UlS5YYVWW49frMRAGcwO+j7DOlpvtdPK0YPQUUz574B4nln1juX9KOjaEZ
YHcZXWkSBlUx8X/6ob0K1CX4L8QiOXscOZjVyiTQ7EGk5VIulCOZZvThV3Zffv8Cw1ig8LmLns4W
gxRnDzV0ZXeySROvZff3n3T1o/WymDV89d9OW5lUtsTDXRYU93hRB7RMZgeRrGHLuPMi4wb9h2Id
KJo3+SDLozEF8mS+4GGbD2Be6A9ewQn2slfsfxvYb96LcQMTx5Kpx5CT+hGr8fnuYOhHE2jZnah5
ZkMVYGNae6Jga3pv+QatfE13dNsMGQPbhMzGyz2iO1CI99msdh3QPSzjIPwYeGSfNoW38GOrHeRv
3iky0h3VU1bmpwGCurjpQfcqbsLQPMDDh5EDUmcj31unoBOcsRofxCytrEIEssioCsgt/qEJmVac
spxbhb6XiSXGDV2tQZNIJ6tKiFiC4NFqhXOE1s0mDErrpo0aCxwcyVZGThXruOU3Zyz8fx7/4J88
S2KCSWfgMWavTIYzY2dLiWa3IOldAoIHA2ucxshjy2J/zwpSwjAdaXPsp94UtcESIYHPnWkZoDiF
RoiTUnwuSEdGmPkxyJUPJol8gzBirAPZC9QEI8LtfIG2lrJnWM7j/pVtwso5GpVGoeSMKG9U6/+x
0msSmDFvUTNmH9MXz0p3fWBEhaqrp1XSeQqkUmACoHKpP6tq531Q2HJE9I/3i1FdArTck8zXRp8S
0eP3FYjFYPSrnkKyEklpF4V2LNR5wEhk3rAcQFeNifcFuPesLXEuVno7oBUgkTD03Ni7/gPuOvVA
msCy6dy1MbmQ0cf7U22VzDh8SSArEX+vOUeViCnpg9y+dokUQ3f3RkAhL2iXyxJmGf3fBeU+0d+j
7+DjOY+HWbPasgOvRrg/FnTvy7zSQICsxweFgtkFJJ8vzkm78m1swE/+sDxXmZQv1WPaaJXpSUiG
VAy8lLGkMPltIDRG1SE4OD2nraOGWqYU1vkhT7azfjLDd/eWGEoQejChr1K1asbvKs14vSLBOsil
BqB3gCZ5XSuUOYqUQyg+ufN23ybjgd7V8n8NtUwDTlcvbnQDj3/OdK6tQqV3xWSozMAhyxVsdzrf
85E/Q1ervBZ8oQVt82TkMGV7sLeod97HGLDXN14f64sZ14mlQut/TAxhCTnxMUpzGfzggI58JZMy
XdUVb6W9KOyWnyFDnUpFJFSdzg2e2LRZA+2CK5TbCeHdLzd4iczrG5zAS3ZF/AyZ2OpizIxxkz7d
6Kuiem4B5iWxDqAPBn4mxWQQTZb/OODT95mHbMnx///ie9lDeHMgjYmXP9Edk7DGyLk+C22DjADf
GAes5rW4hN0PUd8DP4/g1ksVS+Zg/9W4BWtjLdVlQoKvm9tSc+FTk55Tf0FS1tYa00EJ+xpDnOJH
npxKhMRm5+LFYdIq0twpciWUwxC1Jji4GNGfde5ZrX4xGXMGDKdoDtbKM1fdtc4ty6PLLB5K8mtB
c3b52soHOL1/DKGSWyWE0VFHT6Wc7RNOIom3/1iQLPcTSQDYDp8yIC1GA3My3ncpuPefn1bm8mBt
pibaFxw5/EwBpEAHpSeTVBZvIthH82c/ZZqDjS7X5I9c7AEBp7ylcLH3nYMHy7g5ADNexEhpR0TU
EuDtp5j89ntLGuzCEf7DQpEdKVRl/4CqciHakrxq6HFZr8rjpp9s7/0Lr5ZIO8NXIPkS5mx6WgU9
d9+2Nmu/bEwmN2cHrSmIAf0H5GPP4MDLh/zDrp684cq10UYySs/CtXUiTZ484HcU26EE0kJUZtw9
G4Fn5fBYlhGCnowY2S1odNpsSWjDU9duyvkt7tjDTl/o6fVOW940m9Lm2TUDN2qHPj+tPSh2R8VG
jMxBUa4XnP1OOIS2xG7J6tEFZeFIdfTyMIjxDzPLxBh7J6EqoagYKKF8F5xkDcodJyIH3BW+pjiZ
SAUNOgptzE7Gx9/2bbwGt5AUKoyKouQTUMZIwQj4EtZMHC53RmVOUaUdDJOmgiGjjpjuXci6QAfl
t1m9Gx5iNVJ1vk5Oe59uVFdIRJhSVJg8q9IZDuj2qVobVFlG87BkPl7vmeMccIPFgJw/cOy9eSpw
4RGfCoVDZh2Vs0KJ2QysJ4jzwjkMS7pxwuug051q1uI1Z5E4PApwKAU4R0TQT/SvAmrAivJ7Yw0N
eJ5BCT1XF0IhoLk3iSDPXtMZAa1w+Ndj3l37/6wDvjwIuUSgg0nnAIdyxQ86HJMqIOEYEj7hbWqG
j58pPuj5jUcsP2E27r+a3CEO3Vy+MzeTK2noMmxrqAu3PhG0O/+UVqkMep06zgAIsPkyS6lNOS/5
hdsuZWUtQd4OXI2clEJb+fQShPL3rHum/SIBw7rAyIkpbVA0SOy0sqR9odbC6I3Q+5aQdIfPojQq
3gKDW5wZJtvQb8Dpn6rQGXJ5uNyQQjbm8cZFQLbg6UoE7kQkcnASuyjlVe7MJHEzbw2j3wGDITR/
iAaVOJbEViGShPtQ5MyAUa8Qtgow1IygXh11iJuDsgqMaV6YYhvahA4ZyUsnJdgAnG1HJDewyaRV
74c3HDH0BpPnECp8pCwbepRLi9Jk9rx9MkQZUV8M+hr9KZ/4EZE9BqScM2gF+z4/pfDiB/xgqMj2
+4fYgskxiJbrMWSg/G7B3Su9IgqORJHBkb8wx397xeaP95DqD2w/dDC8+oHhnQpB2rl2AoKeD4hA
7Qk1wUrJFrG4S2C1jQ4rRqZejMUuNOsWTfU41k9NuBbKsGI0hvwynZ4tuNcpwJ2OYlULVyp9a4+r
vrXORpZHUmgoFG0g0b4IPTVFlluUlWQOOcKFtCwbQjFqv4JgwD/yCw4zXGPNq2NfdKuO7XQeeg9z
D6fZVA0M0Ud0wMUHn06B3S+i5hkgTne2cvAtLu3JkMtzyPmjO94ahCAxUBHsRjd2qm0RfT1kP7lc
4rCw1Y/phsFi+viSc/l9O4oFsuFYe9tQc5FbfjRRRQHI2b0wQoNjResjAW+xTM/XDJ6AGFym/A3s
XNZy6jY8VYF+H4C5bLam78mb0t9GeT81FcK3nPuhpGQLID4gWoer3al+acSotJM9GyfAHLidcG09
xT6bxxEqX6uGq9bsbEGgsV0uukI1z1mzHzvgTGrXSCh74yYMKx8ur5CluFjBvPDVdGb6LbNElegZ
DN0vgt1JHm42xGN5zt0ooL0qLaFAdU9+YsS+Md+GohvfKPOojcVCDD4qzApTSyBr2mFxsdAhpEin
WM5o1cUtkN7VjAGwLQrXWvPy+tHXOdJOAHdzqbBJhQHJ406jcRc+3+Cdl9x3KI9X0vSQaVLyQYt3
mAv+p4CJ4lqb/FAfGBIVjsgBHCXdTzU4wXizSvD/o/lJt3CGxjxm3kpLxR7I1a74cN88iEpkZ/2s
qK2kO+vKFm4CG1WTNf5ORm+LuFN5wBTtlV9/nEgVSNEVUHzZ6+teZhh6q5ZscO1fxAa7EB0iiwST
iNA2CEqPtBw9SdFCWvLwMyZzG1pq8sxYmdqF1n692CEmREG6WmUdUVsOUdoKgf5ePXlny0llpQZ6
yviph6e7T7+oNGnDp58UEIpdGWpnoZxQa4LoYVXSQw5IapTNS88AjUVF2KBp2F7YBj42QRiNNSd5
B0/5TDTOptFWQ/gbu0WtxIskLlHkw1v1BZ6/Fn5W6veN4tEqyhF35UHZtBvpU8b4xdB0PpjUxwu8
dSFYSPVZv/ENrongYldMAA5+0TP4YUiFkxXuooYHTnU7NA4wBRz41lA21NYLu9oa0z80pjGgUzxO
owb7BRoZ8sida9PImMtz/hcBy6YC6CJIb94cEpOT6rWE8CZRFpxAxJoVPLYk6wBT5NasabQfY9Td
66QK17Xk/2YcnARqBdbNiFL1GC9Ztm8Rj/A9fJtCXAnh++BUJTWaQaOGZj7QdppbzirK4hcEgNJR
WTygQ2AZTVHICVoYlqJU+zD+PQV6KgMJ56TkaHZczCb8oevSpmTs/Y4zAFj4Bh00Twdg+AUq1l5s
gAOF7kXNEOpEVczIaU7ZjUhyimXe9wMXc8ejAGLhK/lwXlBaC9McAf3GT7pr+TJBwHQ8SqFI6M+G
9aFCMqUFCYtQVNV/TG3S5aeYWCsype9rO3l7e1U32b5PgJ1O1CCDlho99IDcwnaGQDQZ2K9qJ2eH
jPGGTWEK+lyNEKvuNFUKbGX9PICTmfgP2h8TTfiLkTbkgt07bELlP6x4G+tFIAMwo+sBZQXDtcnL
7bq1KBWqzQS9uE1D/O0w/L4yFUPQsii1sfzB2mKtE2/T+m6/Pl9YYwz1u3fd7saS0+YvLd38AA5Q
7vvjVDaes4IIi3eR6Eqx3wxvYweF1NjAgR3zAbUGT28nOwGBBqC4bb51kLbzCxWFUHSzeFLbhYzg
oHp44CoEb3W4lMxHRgZz+wj0bGymPTdph6pVZwzc42Slkqy2GABA2t5/g6BIM8PnzbqRJrWpdWmy
rLr0xxo+I+l5hM9ta0kUi4We+uwmms57VW8vpIVmNE/pV7zpfPDNZKBsoZFD8dKOcsUV/tHX3+xU
toEFidYeQuBfHZvFcoMmE0nTaTW/6RH1hlZirERxPMWw+zcMrOTKnl5S0ePC4beHGnAAiG9rdgd0
fjr6c6PVV7Kh7i3yru+MXM5WzSlSuRAbmBLA15y3kkYPZSOu+2iuKPJOwNnLx+RDgTi5cduVKBVk
whvvBsQWkZXsfSDXyBKk6gPoprxfDZGkKbQyfWE8WVmhzhxOa4FbQ1Ijy6uH6lth/FL6FntFs3Ce
zpXkBOMJ6YXXCxFxOzBK4nf5s9GLRgHLPKXa+/BSkAectnLNKGQSQJMnhWMGsaIwCPnDq9GVYJTW
HVfKnuC5XO9cYYhnT8O2CLESRoy1I2OrmIU8+m+G5UD65fJsFBzag1FvFBc4QK1tFW2LOmWqQCay
a5QsvTciq2YRWeBvKGR1Nh5ZB3DwsMFLqFvOqgmnVjwUZB3uDNYVGriwG70ebYRzj1RtqTdOVS1n
3Q+6pqtjtTl6VFI5yhZu7NQkBhoKE/Oza8hU9ocf/Qh90cFEcfERxJArvXU+hUMhQ4yToVU3+dx9
G+TvchYHH0T3LXXnolb0StgK5hU8HbeLIg9sgyA48xYfdAskFvxDqP7HeLI94MyeH4358d8NGU5e
8h96c3xgMsUOKLZcchf82tXXDJKJpLRBXgfCaX/b3x+V4tjpq0FRwcnVyadvxNeBrpbSxjaP6kge
P+JeXTm6b00qC+y5U7a2kVEsF8Mdbpv9Ke/kPUBWflKxud0JRep0nA5Jrv+6TB0VovW/Os7ebLNK
bJ7VimRoPWxN4RtKxo2g6ZfrqvoS9S0H5YMG60wzdrYIBPtDDodAnzg8AcPbszwwfeBvBBd2iACU
Z9Mp3eXwCb0dKHta6RLeqsP/7fcy81KLBNCYaA3ZQoUA9kSZAscUe0DNQ7BEvadeLpSE64us6XFT
dXCyeW2SUNwMcsuMqkhhILCj6tcZVWJ3K04d77URkA4/93kFw9qrRFYcn8xW2zqI+nnhM5GokYuE
sQAMK0d9xEhd37xtYoIdrZ1ptwqtFyfpjRwcBTXpp+6XTsOiYDKPkQ/KA5zwtogBTaUPdEYwnSXV
xzf1Ff3Xblj6dLLu13EiDWKyAzYAOeARQzivrKPFI6v89UnXEpRRNgOaE5gKupiMycH8fkL7Usgo
AxLMwuDLIWphR2eSuiNh1IUoQGVhyaejgo0rEbKAGjBEV7vQ5BSkq9oL0P7gbtzVa+YMQQmVtBjl
KIrpzYrY27ciu769j8jQeiseFjiGQjL/MFqDhldkMasF64sk3O8p6phELOGgAMH017RcJaXekIUW
7R5rUM0lQCcPNE83tQ/+RDzGOJCNUz/uGXIxFBSYko7cgE9Vh1rhplYLysk7lp/ZFgk+kd8HXqac
ExiNTf7dk2q9snKKtv/KVL9wMuURynJ7DkeRJ//BI/86OzPu34yDNgweN1Qbom/nrvSNIynixuww
RsvBtuC2PyfTCCOajk2XREXWjmMxMpkpnOrPhLA54+R/CvyWdYrF5igiggJLO9VSx4wiCjwJ3bg+
PzH8X1ZBYsaXrJiT/ArCblnhitWEiP3hDWtPkCvoQ26+K8rRlbgaqe1Arff0sE+WmP2dSsRGDlcD
YGOX15z/iMVCCvGWvbfSJvY79xGxacrIY9kQ7wlh1S+WfwoRN1mj4ZyeVZHCFWGSC6xhi6qxgvIz
QGtdV5KpVBADj3gWI1WHc0b9lrWdMrx2LkqVI+yU/XDiQw1DUpChTJEMPCiFaHuL7/nSopNXFt4J
GmW6I901k1XdCy0yVJ8Q38wDka7Y8HLC8R9KqLiBPuWDHFrU+5vZtAV3KEN/6FxhlWoSQZESMTid
E8WaMajF0lZpjcbmRW0reAD50TRle7Wh5tsrCkVbwszmln70Nn2TPv0izAX05MReRPigNb0xAEvv
JVumK8Vkmx8VaBr0+Mcu6THMB56tVlgvtK9Ox+tq7fWLIY8Pmje1VeZLE/8ejRK5+a1+OZVded1P
HvBL8C9/vRXbrJErIOBb8xhLt8oOVJ+CqpWn8HQb2o3SdE9qECjNhFT12Ct8V/J9FosLhQq3itq1
RVTCjSpc0iwjOXuzi8GY3/n4lcm2V5ByPomuDwqarB9onIiDcBuepwHa2RlS56Io2Qko826f0FB9
ToduUM2YNhd7CJS2Ex+9ADtRMDPiaZAdnhibDwtj9xufBs7sWs2srbs3sCp345qLf/rejh+VNfZG
pP4S/VOLT1afkyrmdpklrO4nqw9qUf4+BQPYwXlaCTA6thkd2XW9T+JZ86fje/hWZpBdU0QES9cv
GVsw5BPJowyi/Owq82X04JawGqk5Lom6NedLeCr/a6hkGJ7RNXjXrG00mL0qGBibzYUjrprhODCQ
jVDx2pgy7hiMwph3Wb69N/xBdd8q9l3otbX8nkjFJRfxi7huJi5gvCd+XDTT0NtA+QSUdJlyBlyh
UHfBjmG3vVWEQpolyQ2fUPqV0cPlfdUi3TKHOzyTb5Sgtl05P1ksDM7b2aBG8mQtgdVp4hzMQdzU
Nl6ru1896pYZu6AfLtGOltHYi4gVdMNWeKRkBslCWIm96Qtw6++fd6yFvz2SB5e9yZwsDCUFWEwR
WhB+QHL1ODJDbX74RmqxPATIKjO1liE9eqKFBl3Ec+shFHk8H/QjxMOxSgc6/JV7cLFMX6IEyi/+
pzm7JC0MnSSC+oC8lMNNMToW1Zqmi73Ew66BfUjqflGIgZzpWHZSCkXjs91l+BM2tbrUptyoeqcR
n2ph3VCZe6+r/ctmQEe2mYaJFd+9PyxNslEvlKiajUVk69y7XWZkjiwwo1b9ZktRWyGO27qFdSTg
jwVQ2nu7zboQZRlZqO7mxm4KVKcEPHro/NgVL/aocK8vdC6wvGlK986oCUUjliQD3drSb7QvE+4i
NSqcEq+Uvic2YN1m7IkUE4w7O5wYsuU3tIApzg1zmPKgDBfMxG7lnXYedBaIEIhUbVATLxAnRmLn
MsTtjNH7Sn3SlJqDzVLRzPh7aZMOuvbxgHzgHF5qETk6zBMXxsMJ2q7A5b3afFcJ+E0QyAmV5UiD
aBU7zD0wQPkaCnxQ/3VV+01wmDkvfhUHx4E5c0EXzRw1SKhSbsmSPHWEjV8TJH8lbbTzhDdgHupx
li4ond6iX/l8A7L/Ze7uyS1vq+R3eHZ4kt05I4JN81lIpOhdsoZFM8UeVPcUcpeKsAnoBzbsfoBK
tSWNClTmDdSzR820F/wzPsBlsM3yvbyrLUU/iv13qUZEoRIgBkdERUn6UfdH0P85nsz7p4o2Akys
adCCoJwy9Gxv6bJ9e0pyeSrEmeRSbGglUJgCAoPjt0t4KOH6mvg3t8xW6FXslmbPSZZ9HkBZ5gYs
qY2nKTrNf4Npivr8B9E/mggv7Itbc0zR2JyqxOmv/seUJKlJte4bP3fQW6oD7an7TWKZMRMMxgMR
+dE8SoiqzchGyTQ5B53JmLPqChyx3LtF/06qIuTTNZxTlCJOPHZKXZ0/yrdHguy35zdW3s7nDbz7
ZInphY6rAVTf9D9crfyYUfE/jjYMcg6Weu3D42mz+85NweAhwJYpyAZq1rhjkUQZjVt2IK4C5/SG
NL5yAaMUEEE6VEmSiJVa8Nt6tH9vTQcX+55GLQHAX1CjspXAFaefYtY89B9XVJRtdl7TdVNEZu//
4eiu4fnCRgU8bVbkX/EwYh1JP6n9z0pyBf0ILBDF4jXLKbkNtO5GnIRCMXTmnp9FhT7db+SCsju9
ZvwCWC4V9VxSwU2FzE/ahnz7NtwkfEGXJN+0o8CwLUjGVBrxhPetikQp4p7Vnot/GNlaaC16TeJj
pa6oW1UO71yz744/tDck5UnUFFabpXwkfm0lGb2lTSAkOrd5kRxXVfhHMNFBc6IpmN6Yn9/P8QoQ
R/d8w373ijCeyhwo6U46gAblxMkKNnG8vFijdAse/1tbiHxWgVCEH6kmSERYN7KoBm99BMEtpybi
bgvCDqG+3QGUGbQi3LyL8A6ob6ZH40mOwhkRNToJ5gs5Vt0eqryr4be0ZoJtB2O6SMy9VtChKMsX
elezc+88NE4CZDwppqhTZIxBPGVisAKFr7PMOmjBZsNkfoG8NsMJBl06IcqgAnJlCLIKwJV0ANyl
95dceSdwMhLAz7F8TMKsYJxhvpxt7sTYg8g4o62cmkUFxEslcOQTB7yjQXpLRlAkw7WsnKgdlfCb
DaXfLqAGhIf5ixuz0S9cYcrOUPf8+i95u7dwW18g1Ti+8MlknaBvkQF02nevINelSNBfOwxmfIVe
9JF4fEoykaQ0vjS7zs9qR5byle7lvTFOextktsfGe30p+NyiXTgWTXoX0pU6edZ4x9aXUnrT7ZFj
ZBmEcWgodAFRYQijybaiKxA9tQJXPPY5GnY6R60OEIKx041/vCApZvTjAysQhSU0c+yEYnR39WXa
QHPi4jHPZMvcyTnm+koR/VS3hLHK8XJCHAjlRwhpGz7+9942MjhHsvYa+TWUpyy1c81coBOWY3ic
fL5cCkba4GXf7vLb3/rfcgi5IbpFjXAW4rMhoMKqfZcfAiAhThO+7TFtiAIgU0xQdLVWanDd5MXV
0+evgdeV9HkYjbGwmMYxH9JPNZEch4EZChtM/vs5ERU9i53D+3Ae9U4AmODIsZVqOcCShLlU2cU3
hOAFenmod53+7mgVcg1yLzMKPcdtH4v3pSDLzTWvh7yVjetHwFwjOlIVdSDjup10WlAmNxasQEq0
SCjMqOIsD0MWgF3fKVxN5ejhx6jyfLs7ETA4YIe5Mjz+1yX50n/FJ+z2kPj7Jomkr1qf+g9j+Qxu
Veif9/5D23vk/RB9Tjgmx7v9qWhiDfY81ELTyAq8JllZYqe3XNgXaRYJZF2n1WO2fOTERbN+1Qy2
hdu+6F8YjTTQbIQ09zGlUVvInQmyxLkyhpNAf8TlW49SA5p4Appdj8bDAvKPdCumEssqMwOaOi43
Sviy3qWsZUumvrDz0HvUFnVOAABRMnFqS5AOcUEutqkmOSzykdDL5jdzRzxCWgYYrzcMFbI2q5vU
+QflvRvTHK5CYd+0eOeZ0bEEXyXJbPwDM4dPkGtj8+iRy3pTxtgUBamhrvxCe8GtG7/UJ4LqxPcE
hjq3pSLZk8/rm6FVdB/chlrWFalon4IWXUsDol+ODJeTWUWUNR+bYHMVVmrPN6kkjdewRMIaXJ5I
W5M1Xy89J7z8kYRB5sBdMbHvyvcONRnz+aqiYnvwdDVoUBWc5/Kfx95xRZz5dohzRjRD1NcxGfFe
MljG+CzHGU2ML9A9d1JB60vTYKGg5lED48PAX0U+4uCyt8ZeZoz4bInW/blzAHD0nno6lCvoEQJ2
937wKjYjKy7mr6FD0XIHtJKQkj0+KHup8OXSy3OX2DedNwZfMGmAGnk8u78fLau1zYodVa+RtnwO
L+yrCWmshDoTSsOVH0JLSJy2SkK/eW8hLC4piqx1tHKcZ8fiaQ6WuGvH+ykRYYJqCMOZiTiC1LQg
FFrNyzfgvEWDKjGba7DvE/COS5iZBUtga2j5SdmJXgIw8MszzEqSxsmr+nB1ApCso3H1Rfd0T/rp
1HGH2dzGcLpxYwWQsJS3TgCHlRzrbYpdLpg6uo9XegH0nPybvdt4JmYFGfcwc3EtNlrMpAiKgxtL
4gYnRZmXQFtYAugb6nD0IXHh2wJZeq66tK8rJpwvuTs04tXJsFjeKK5vWzD65cSfBdGY/IKUOkRW
IdXobjYwDUNW2E/NRoU1d46PGeaHRFjPT3njXHzSeXUnmOVOCvV2DmQ33XxQcMCjrcCfOXkWaSFn
NESakYawkpjtifATiD5x2bTGDD0zK3v4cV8ORB2C9ofqMAzjqhd/Iw4odyoNZo0DyBMExUBbvwCN
dOhEjwtS/hiwpdNswpBUPpauilmKFmmZ5igKCmWmAnd9EvHz2hRpF7IXPeDEthKRBZzjc8jXuSJ/
9Pn3Hy8c9gSUhvz1VS46o147hsZo1H9QYf2C50QCjyA65mflPYZA/LLLNgPd7C/ZMwvpMjAwUMN1
mJxVSFZoRdVZ4NtSeqZ2qCCo32YhaCWsGVwpImece7MDt3psBjunVsDGSWI1Ak9RzGsv820FhIdM
BtZNc+nArMUpSCVRTlDAfFf+A3NeyDyD7jni7nACEXgRVBuNfMXMuDff5cZgz66C1lInLsFqCjQa
PDdkurJVvTUGMOzRKGRoTBWKn77xEGWPlbQuyhsKAZMR7JCIOcMUJ6gLEXao6IjK++2qhPg2F0g3
C20hfOvEKpCb8Tbo8JAlZAdeX21MDNUfqdAALO5yyQnGZPZY7FyxXUB9EKF8Y3lLbzpAy5/GXYpP
NkyVeF/YO0laXlk//gkUppXOmD5gr/bEfdbXjDN4TKSYv8PLSHBdb/ihJ00HzW6ACD4jpfEkpvBA
2tHjCl2ic/d3IRAG9FMHDN58+XXbfg6SP2KJ7smsO3Jm9NrCJinby6JhqxaD07IeuKztuWyt42mG
udCbZcxoXzl0JgACatgWBp/epTG4u8UyWwwq5EPuulyaieMrBUQ3fjmgoO3VMibYV24we8ijMU00
gyt7DWTGoymxqnhMs3VnLQS6rh//tK5ROLI13DhRXtsgZJeswNCf9Me0D8lemU8nEwNUBnQlxkW4
lX9Pk10jQiH5L5rrljNB3RYxMDmXPzFHS/wAkxBKoRQHAgQqfvqaX1QZF566GYoZoaWqjR6O9vb6
ELBja4NikvzwbLyB2Av+fPSzdWxEdqLilRMGzPcSLIcn4g4h4OivNI8frz03TdQMWyUfhzVzo4mi
b+n+yU6yot5LvCb0/vlBKaW0l+QHEPMDi6dlCT0O018Il50tDIYiFhnCeJLQamvZfbbLtopk8im3
7pWwNEuGMZmcmjWXMof2MAHXvZRXrmuUNIfbFe7RrmbGn2O4K6Yx0rxVEODmzgIfVL/gt6rqb73i
d5NUlhy/qTSHsJvrb5kHOPzzN4EqN2BAKQ0GSywWqRwXrRMW8kEx5p+/MMTaU691se15DZFJXV+A
3pVjyG0UkebsrJpYo+DBkBPULLLgvMf6VuJQ+vgZuusLX7m1u8yjSg9kR+nCgRm0Eo0oRVI0tVpp
W43cLT5pmsItYRkdPgBvpw8T4iYh2faZ+/5REFr8oWj43Z8ErSadtlWkI7BSg2hNQB8+A/FsWlCu
rt3S0gipRJQC/UFImzL1X1ivYYq/hXORRJ3siGmTPeb6jyLHUV5AZ+SDRa01vLqeEfVJtorTCP1j
1AcEyIKHSK3eIo7L9fTUO5B8bVaO9kSibxhIyXrImArhLBpJCk0KfflmD3Qj+uQ6t6BSDqiZBoHC
FUz1P/KB9pgFgywJUunD+EROSP5EeeO86Kmo8YE4thaBibGagnO3zhDm0uQbmbU3H5lKVdFJ2HkF
NWBJuV43SrQbZr2HhzePr5LS2Jo04qx6CbBXbI90xaEMhEbzm5ovF38wy6ed3cdtzxheJTwsG4k9
PXhYVHsqBZCuVcPb74N3kO4TtgIwxtQUhXpI3puOQu7DixDAzFJbiEIz0mZORkcKB1KoSHMD+Ofg
+DIBAA7+iNbyVbuiaL/U7wHh8ez/6PrONtsa3O007gz4A5iXvT8tqNfkcJuGxg5wBoEUYLv6VR1B
SZ57MRoSn55dhZNX6FHeISrQ3fxfG6EQvnju6TksmUGZHP8oYyB37fBZ0f+0h5OKepLOjLAXuOOO
MJzHAaVUyvhlnsdDT4b70FsrhcxkgkBeSFg1cT5Otj417YSagkpJ9RyF+GeakAsm+1dBwstQVwST
R6lZj7AsS2toB6g30zeC2saXd/BMcCV/WiDTGgdOTZfMxj34GbHtB1bSGqIND5MVS1bRMtJQpmUB
eA3Cf/9WjkijSHe5PSZiYB34kmJo16tYOHM7QCEK0IzOD1FQqBxNwQqeiHUUh5kCUE1Y3YzmtDi5
ypBSYwP5jmcOL6lyTk8V6vTw9l0f41hf0SkekPiOcWpo6iyUqvfl7aP3uxiflSjFYbs/j0UAcWQA
3VWRAKJYrpD+AbmXfkRBM8Khj+LH0nUHi8aaJ5yO7HC8bPfinQh+9TJ+TTIyq8tQwcHqcBZTXcqi
unODF9YFWmw4AvEx0F4ObxXp+1VRc1JKwJUJfP6DgfDUSBa1ZDp4B7mBILB7uVRbzctJi8iHz572
rCfDDNwtH6yWyIyoRTXSkV9M5DcikR7eS4WYpzsi0zF2dco4mqZ+zeLkMzxI+5FWLs4nKxoHihzp
htyhUwKJuiSP9aATTDB0Jd2EOMzSwQACWZ6vsWy9aG5lUgEqu4uMC8Ttm7JpoU1rMqK+JaMIBNRO
EdkYlujALWCu0/R85jlc+TqUwHQlYgLIVWW8vnVIbeRMzOnBE7RqiMf5l0tV99NQZDptyphMe3fm
APd8dO+HD/HYQV2uArS3vbLBzCypYdyFQmE0LErCcer7oeJDWuAmQY9sBsHsum1PBw0ETy0aYp3+
/6oIWG0SQkajnOI76PBgOChXh80Y8KRVOiyMYbAKbpkFel9MKHXDT2K+V0fh5IANZ+vmmMDogFE+
+8u0PmeCCJquNEJyefTyZtgWMUyw0PUUwINF96OnjtOLVHcCtC2S1xjjkng7Z8LQmmKOudL8FDAg
PDxu2pXbjss5iyqZqvAfMT/ut7xa2LR0c77V9cfCn/q9Gd2yYDdwPXWLv1WGQwJJMhybNvLfZpjJ
A8RHiE8Wxen1/X7vs2DR6RIM18CR5mdiuBdXZhaT04r8J38fYFpom7MTirNe/Ghv7G9RnDUOkZ9K
B2cecxHcswZ5ndP68V7ltVOVF6dyxNw3FtjLunOBQLiYc9/rHjh9FntFgAbyimN/MVjzj1k5T6DZ
aq7kkFWR5L8o6uMvSlYDJXDnTpMjJkWZmap6FcJwYwmthc9bv7M/10wyPwvMSDN75V2MO3uo1CIW
kXNlL9aAbJDI8CoZj1waqceXACX+DnYCmLRF7oCXgGQFMtLP/JVXJ5v10NDzN9X/bs+6tKosq6Cz
3IJT9uSXjiqIU98AfP7OX90h/tr2DJrdtpdgD6OrBjgY+5qe+t0qfxZujqmRIJnrCspmP7NkpjGg
CHoOFCNQ8tQyU2n1zbRzn+uvTXVuMgVJb0HtQGvAru4FNK1sqV4wc6075z/vl0ayuWUnmjK3M32P
KOxHietFVdK3aGO8L0Dk2YIeAGk0kus/6P/j3mSgi3rcv3pvHv3mPdyheYF6UiI+T0MiUTax2eqH
ygyHpDSZdxHsqzBrS4U5cE9Nx/Y3+t23t3KProO6Fz16HnXNCx3nkIBU3lsOOY+2qShnMNx2hscB
Yxf9np8uNPG9yyqhrBR4s1GB2r4eJRuSAD2dEw561YZaDjZMdGoZUryLPOzO48tpCyBKIcR7q6AN
F2LYYivhwBVjReCRoOrCwfC+FOGwN7Ph0CYQTjBPO//82WelHzReW34EI56qoawnHIu/ssSfQ/Hg
qqpZxaSps0FSDaEHh22CBtzgE3S54Zznm4KfaaY6lD1H52JdC4+nj/0mRKuVqOfKGyPNmqQ8b9IL
nYvH5YEXwaHoVfbAcEc6YSxC0/J2ULDD6zt4gojrfPe7ulqgeJvWzUyH1/UKjYSRHRAFYFOwnsKQ
IgOZTs57jA5PeIOWGxEOutfaRmPmilbvHuLFekgB2MH3vgDMElR1AkLT63a1ucpA6TGimpVzOFhG
gHz4xHZYwptOaurq3ft6Kb/u/dXXl/9EEygljWRevIAp3AvRlmvaSWBYGo+gTnPT+ymTv1/UzrkR
EC5KYJApLuJjDTJKB5io3cSl1jjaDq/TRNMTwB6gcB7jKLqYnXSpPWp+mVx/p7cHTytfUOxNN6if
zOlHWhzpzKv8WbNgjMuCZOSvOk8/VA1c7QK1sZm8SQ2+eEPiRmnFsTUxeAz84e7LXY7baHYAJOng
msr1fyB+JQVrj101rVHEIjraQMxhnJLyZRRJkBvAZOPEE40txsDbTR2NUiUtRIaWciN8iXKik38G
KDjWnFCKF74btI4QDTFxpnBPcdutSCOrSS53+o+HdeggAkv228eJe38yXQcD9wktxN1GglZrocu5
h5MHHzYqdHW0Hdlb9/CIjwzd7vpPJRkGoVGQ/Ak81GFRn+rEj/LTALbkLbzxbWV6uMtZosdqQyMG
tqd3rWpzvLnYdA6xdbWsFpW+N4ARYWvXCpDUa1EqHrA6XJ71C/x5fB2vsMuRqipfnYEsMOc0Uobw
6YJI5U1u4xeWDk2aYoh7Wr25Y6bW9xGcENJOluVs76RVk/9/oppe/zh8ZqIWbk48D+TsUj/DhmMK
HgUOwD1RXHcQJIO0mUNjfbvLXYzvp+KhmxUFftlfQoYN005pF6GsCGIiJbP40lJ66r3RFa9pFA2r
PschpdenIFKqxDYB0V2xADtBGouIhiM3EYt4DMblOq4hY169AzVID6spm1jVX8cS2wsHz/bHvskI
UCtL2ZLHUNNrV+5+0Ze9i1cpg3fgnGZfCRw1cmLyT2rKsyB/mpr9pUSH95MPKnknrc1QO9TxPt3L
yck9RAKe0k8cjYDv5Hf9stuuEyewB+TVbOWUk8lG2xEjVNhGwoC3WbwHy/S1B0Ie/VjTaw/zaw2l
wA1CHNmOxKhFvXndwqeWjHv6lwgyRzSy3PyCCk1vwyWsTrkAiYKvbdUTiRuvh1HuH7xNuG6ZokEf
CE1xnRa5jlK9Hz73bl91JPeXtMNZsM0XXa6OsFXMdaiMkz/ANn68K+E9lgIpGeHCjCkAz2VukZd+
REtxI+eIDppRr8JCsfVV5y5ycZpgW9JNZEfEXtuts2o21ftz9g3UvX0FAwT0I4CdMZnAl1CYQYov
5CI5NQXsLAr2x+PAc9A+51+SpFdWzLIWeFxvL40bNXPYCAMCGXff9P0lh+Qm5FvD8+tXblXzTBPy
xwweiDj9OLH91ZEmEVCwlrGY8kAg8jO8iowNnw6p0LM1vJjOrf8ZmfcHz2MYVS9M+xYZJUfyK26+
sE5hYo4uKhTU3u8QUI5z5K55zOdhzqt7iIgksSI3HypxGeaf7X+iSX2eg2YwYa8a9h/MMhkAl20W
qLArPMobQu5q77xk0qT9euxpx3WgNvwqmomuYDJAnMlqCu0VBDxyNsJ34pOEiVZqEaYSVvRVo+ML
/HeCLVeVjnX3UORlJp74AcdCCoaYBL5GJFe2Ak55u1P31yhTuOEzWnJjGUoRd7kKIdlXHEYIcRA/
rZVb4pLj++Wu6Ukes4t+kNU9/jurP1XqX3p9pLIvgbH5/V3llUUHCNzLO8xEZZf2/a6fy1wPtGuB
9MNegcSY3rQa1Ky5DuF1Wg95g2VPVgonM1j1z2TaBTrFpHuc3WX6YX2GXfX6RzaMFGoLvXYbl6FI
AMFQFwoucSXJhpCKLkHqHXM0UHqw+sD2h2TcjFtlSoUUYKuK/cVrN9xCA62/AvJJUrKZlfzQDJlx
3hKrYGM8qsV8S1s4JrJZtesEk0qV/4Ll01YCUIW7dK0WWd/EKOT+e6RSKrtTdbat+2LUEBzKFHWO
w8mMDzHxRaCoRoQ5IIVUFOXsN0cEPX3xU3f4/ikt69+HiYDh/ntrZ4GNBjl+Yql36XONqB1FlLOw
bjOdARxKtdBRgmtcvsq9toDl4D/HDhZrBG7Jp4mhRa0VuPqvTrJAxBSqgnnQwApTbMDHKfsvDUni
EAISJyhWpzG2wictGhezfXoyTI9SFqADAYUXQrstxVYdP9yfkzhllAG7sG6xv9fd/1QAWvlC+tsA
BfccH0uDUFtIRo1oaE8qQA1pQPvpZOAQ9N+MPFQIs+tBIgM/JYjuCTLfmCho38AN/z1UIxoFrxCY
1kHDbDvSuWqDmXHPnFPeiSSaCbGwYqmcOMYqQy1iNpwfBPAVwK0XkMjYjrpAHfafQnnW6G0e1DdW
3rEoaJus/zRaufNhJgYIlq70Oy8kcTZMRDMCoYnd9O+KMsIR8QEhMKe+iP3RmmNzjGPaiOyNEyNP
uxNqcRRL+SvUBWrwiwsjO9SOoioDhePNkcvhK9ZSdwq+MOeE8pCg5kG7aXYBU9+/G0ZnzH6OLcWc
ynipnmQqQXWoV5kbvXKiVkBdu4wnhgf1IcaVmg+M+LFc6hJJPrPZwU7kK6UqIYHbkwrz6eW3dQjA
vYyJAgvLtOKdIqkM5Npupm8SPEIO8tvmEgoON0AcLhRzePBZWlicaqFrAfxUCa5q0saZnF4MMqDg
Jthqx/GdkrVsVtqo/O4Jl00ONs4n2fFyLI07LMHvjaqwQuYUJjl+SUtYQ3+BJjuQcjaXisPfcA5A
eqwYfzucGDbsx+yzmQWobF5+Ea2y4n5juLiunn/up5hNehFTR2u8RzMQA7s1D9QzKtZvc5IBl4jn
gcoCZQgAiX2PcOT+/Aoun8H2ea/5wGUYHKgojMqnf+qGo8rpBxQ7iXpzYCNpSl3+U/noJCAp/asO
fg0WIxdI7NDsEmpMv4BNLIvZJFCloO3YvvwpWHiscrQGeYxVe/m+8fjWlL3aR6HVQcwqcpbQL4Qq
Ha2mQ1/6yQnVOCeWf++/sTo4p5yl0CysgS5PfdZ5yChls4NWGICq8e2qxzRUph1X9S05He9qJVNE
7fe0HNAl0sMjo07NPodyYjuW58sRPQtqld3eTr2AGu28tcjOy6eTy4fly5mprJbGcDSw/7xurEZx
IX2EKfmj2dZEEfp5NfZrAQbWjQ4QQpda1p4OBZA61r2ihrRQWWCOKDISnXzfdTYys5Nucq6zK8xd
y2I1L2Km+NSI6jadVuAe+lUOougPv+1vFbqT3zreSazuCHHqBRcuKZRAsc0lD2c9lMd7rg/hYYBx
ppvpfxPQbeeGaSnHgZmZCWK0NkQRNR8HuDvm/Aogb4m9X2iurMjpGslnP2+pjI5oTkW9hKqh2QS/
1wnFG8IOPL+JPMPG6/iQMHNF2e+HvhC3NQrIGSAngbuPUdKLjO2Hukop21PO6o3JP8Y/1nrS2yK7
okVI2cSNccXix2qP36GAnuoPenzRcOW/qD/tAdU0w1NqlbapkCknhUfcgzkIxA0Z3H7WjPosIOem
7AP5KQE+glW3UGQK2i1pu5v+jzQ2J3WVRLLjaQMCHPhw6umqEPqdCC1l+7TxV6mYIC3AYw8Xzy8c
wQETp/LtxcAlQjS5s5rZsuxnhKV/kXzpAPzGZZqirf0WVrfK42AFFrpsBsm5TzEIz8lMvt0M+iqG
pSiV9X4FQcxx5vFcAGYkQ/aEN1D3Z62Be4tsJJEtVsibct7XSWPDb433b9hhjW0Y9HCBssm54iBM
IflGtM76bCJbRpxPYCN4WjTk5xvwS2PWBoSuvfh91wYD2tIJ2yI3V7KU7DkiQwgePb78nM02ZscF
/Z/m5ei5FiaDRCUvpHSOO+313MFIn5OTjECgIuIOMFhXFvzKpMNdI8eEn0IrA9CiC3qnu/kNwN+B
NOIsMUrPbR0NjyAwpIJCB4+9rKW1RZsubOEB2LVqL6rDR2zRhMcCPuLcm5bh8TZX6ZvmaQyxquON
PXh7t8U9t80CavuY1Ndj0W5BMLRvBKE4PG8OezdHsZeg/NxwNi/v+opu2Z3pNc9h4Dd7T+7tuhKi
AP0DpkVnrSkPUmkRSCJ1/OuiFdeIUdMRmx2JNx0carYuSpq7vlTby7tV0n6FYi69z+BUZDw/7CvV
6/QeCujcpgzfhlbJ3GbtcB9xy74KcxCUZX+Z0ZQlP53FlJDW1dwM3jpAIIA8LO8ilKJKhCg6L1Eo
jQIR8wsxym+SXMkVKwm0OyezEJ3ADhBrOeFgnrXTWLWPQerHh9l8GeT7l7eL2rXWnx6XBnfhPs/1
pn+mw7tvmfVyybFU4ihLMk6rMc4dytyomczb/nymtRiMnkar66x5dQe/qsJai0ab1MWI0tBmXMeS
1/ilUHB4VmSZxZID/mXeoxkofebXHdHRdPTLxQ10kXd7AUtTvb93X+5eBhG8e5adglCxnhYGwUOO
HFz6p9PEPr0vZOv4mNVjd1+36Z3RE3bbrQTq+LdEOYHyFjL7VRwfNBzKEB0tDtsb8VfqLiNuO4sM
0HwPbIfcuQJjvQ61QyteDDLIfso0/OBiczBr9oUlkUuuBkoYXdK3h8Ud1Buv8mrLPAtyIKpaF/wa
kFDWI6kmEBJPugpGM+GTybQB9wodpeR65dXsZxXNNCKWEXdP99MLU/tqqnI8CX20ePSLtvz+8Wwc
Jcz4WjmtRnM1Yx5pM45UqtwOJgI+Pr6o7f0WxfGrJGIkKRIU0Iej3Lovzdjsy2u9DJO5lR85iRjm
HLqwSIJyBwLQVH80EFIwNfMYzjjNJwJG6O01hBeJix30jwnrshd/RtIJnVv/k4K8c0yEB9wPCMxD
RKKxmOMZ3kzDkv/tH2ZymblzPCE0275c0AGmJ9784g+0PiDx9gs37pDzY4dwTDpRIXSQHU/36QYm
yusghgu4989W6oXd6r6VpbaSg/7CVhit56/jcJ2AWoTuu8ksEHmzIgURDT8K6hzjS1iu9cXK4ukB
g5nscHurM9HHCA+RY4+4QT/Lwz5YS8Cri19Ukt0btYTljCeDmgkIDaTe3COMiNbPbQnv1L9+6ELL
M54MOTJCZBtdnPT2UOzqI3m5bMzrd2B6DcNQyvnxQOeFjhIqBJiD2GZ6tLW9v5/O4uTxesKFoPki
A3lqLelYF+ubtqpb1vpaQPdygMj3H8qTN9+wkIX5/nbRzuywYq5Bp9WA9Ue3MpfzVfIYcwW9PXLI
TqL7/ndhov3paiJNqBH86shp5ExQWTfJtzSgQbYjsuUFy40rgRKiH1J+rNLBd6/Fukqca/TfD/c4
2hWkisXACTseJzjDwXJYWRlQfS0SSm0mr4+xqBoAF6tHmZ6m4Fg2sZStJSAwcLD559kgZqXrjtBS
L9us+qTfN6KS0IZwH+0Eh9oO9zi84m/wUkwyxMqFJpGm1OI6JX+JQZJrbXNfpYiAx15VVR96lfJV
7LEwvY2A4uKpI6CA6Q8ZmqX2OBOD9xhcyD7Cxd4J3QDECsJHupI+/40UAwN5B2k0muducaHHrDEz
41xYasUd9tZGtPWoOvShRMb0y4f8vC/z2N0Kzl9AHYPwfT2yfXyo5GQd0f6a4wXNOCbl0Eevnw8P
niwpUcxiIv7XxinLhcoJ5Wus0rUcNOIyT+EJe79VHcOiIQvGkladLzX0UhDFMQ9fhy5k2zH9yFjo
GXD933TX6qHeO5rnUhYB2slYNIi6UJNRHGwE96slRQrS/4oWGpDwq3Um/DrzSeBbjF9dQdQcedpr
1qB1ftG0XmhEqNUhlYzCDsUgsjVlfSFGLiRz4U5qFH6scsreRsKwfKE8s8VsFHiuL04xwrPTOJrS
OjBgxGqVZ3d/t5uxa1aLXw1fOM17/eMQvLYXCufwyhGd+dvD9NocL1DDu5aZR5BYxP/Hz370iU+b
v8nm/jVkBS6eBONrjQj6DTHu/dJ2lMfwKnohyj5zyFaGc1okC+7Y/ThC6r47fRbKeovsOnBIaGAG
/os6mT9bxAsgkQ8RZY7O1DHUHVCbVzvXI7cri508EmyQ+n1DAeZSAWUN2QDzx13v94HE86zcCiQa
fvP8wco2kcrSz4aTH/JU8dS6JQ+g2Nhf6O+YwAXi0dfPJ6l7VEEvFRtk55FLoWh2Yci9qPoSSjtz
h01dQ2L/atUH+jKwN70DwqoBNO4aPlpFFZwVG0hkWdNpd6cGNLTMWBvvJghB+BLJFuu/q2I58wh1
mTwq1u3kyrTRfpmK5XKFTA/zRcqNXtGqgI/K0ctxmK/GZskNk4r09CunXCp/Q3EmF7x3BFDkH6G/
cW8QZncUEO18iXXeRoLwNPudqRTTEf4QX5u7jzIwd5sfmEajjg00jZC8LzdYy3un+LG8m63Milir
hRm5s4nWD7yv9d1SlX2kKNJ8IoMwvDWK4V9iq3PnyzYSewiyMO20XcVhpiygO7H2GvhjPxCGJNXm
xMg8CbTKdvl6i5a1br3bcY3v7RkZxAMDrjpPtycTaaQGpMTl30niZxB8AS9zRFqBvPRlibHI238n
bK/QKty8TNehwIshJHlXVW7BBvMZz7hv64IPcYWuy0ZPkUs+rlxOrsCWLfKcMXdvyxLa5yj5DRuI
cWRNNPayOHLTtIaI+qpirFJYPAVePYuNIDwCfH/DKu84aeSTU0qu0AvR89xYYD2Xoek6DirsM82a
+jxiBwaV+A1Ln74gfxPP0nWD/lxxAlI/L0FAkoURUMFp34znJwx2px0X/H5q3HhwX8KPXTfAPEt5
ql2VL4CVDXn5UqSao8sCBXjgdG9cBRfVdT964xVK2oQ+rZScxQxjJPnB5XVGwA35P+OaKIv/J6sZ
YZXCEqenVDy6muIi2IeIfSjNnoFImQ3PdzLCpggUQ9Cmvp+nRqkcnTObVKTaOIRg6letVW4EFg7S
QH+3U4Lz3wfZzQcMKLOVTQCslYE5i4HtDggrRIrjBMWo98FRPnTKTS+88GRfh3oG0SdzJ3XcFnte
y+v7Gbl0BozXWfAUXI8YVRTJIxZbIMNvOwyBZAUGdZ5SbHgesdkkfkC+2sauiHBHPYyBiSf/QLDO
ckS/3lLT6YA3CrkGNIcz0vMKiYXtDa5tB0FqTG5xiZAmZn86LfZ5ckj9ZiiDPU8wBmfFV2eM+9zJ
jUFjzLzGB6ksVwyG62n7749PwsOenmvd1hkKB/CGccHM1mBk2/gekZ9QQ1Fs9GYbjEx3LVOHu5aG
v1YoK1WtI31pH10yzKaQGHBLYV/wQK2oEnxLvb9nLg4fRMqjI9wbX2pv7CzOcqkqG6/JQ6V3nyvm
Mmw+4fDFpc+w52HRMY7rYsqz2obpWLqWwIstrIC+IXIK+sxBCvvioYYNHdGc7yeYQNj2O0I4t9g3
OwviuGNIPNTLGdEkYd3kZLBP2ABKyrjoC4yOsaahGp19tRVQINlSoKkzeUtSiVgRWD7mRGMRvMlz
6MV8oJWWCQShle8IgWS5Y+vWN0T2rgdE3dg+NmR7a14/MGx7ttlgoI5G0CrcBb0Cy9f9PEhVEW6K
j2t1QboFD03sKcfw+9Rv3w6sa1I0SrcJNsrb4MzzxHB79DojZ1LIL/b5xFc6IbJ8tSIdkrLTC31g
rVE4CiXQPPfvaU64JZzdvzWRWxj8nzFIy+yw9N5OP8qbmjjSUqA8OzM08fnVu2dqs9ADaMPN9g8E
81Xp+93RpNE7kCa+F7K/JDwQrhyh7HI30pjGu2NvVyAQ0E8Y5b34qrPvAAFupH2ZUGAey8AiC/qn
w1RxH33E51Tit9evS+kuxX1GE6JqhYq/spj7t2ChV1qVXEvN9DYod+U1+/VIJ770Ro4R4L5aLpIS
nJLF++JoU+9T70Mvy3MnYOX0RjNx/Pe+iqC3yCLfPaEntvDGZFIbwFDYQqBmlaoFIcfGp7vk3L99
TXmE4YEFwFExfFaq4Dih4biSs4q3BNqGU08IScF4A6UaPhysVG6CG2AKnOkUj9NQvy3UEp2CNm7D
tBu8NsjVOSfhYyzPvu21lXseecIN2UeWQhn6ApOPuciRlNx1jUyfXdWp4U8qXOvgfcUYWU+xgoUV
qp/KPq7teEs1xZFN1VVNXc5Qz/M2vVWeq10Ha8Q9Arg1b7BlvCJGGXcMZKMnGQVDCGsiqxyFmPJt
6/LLXXG/tAjGuO/n9rIsEzUNP/twMSUUyfNQDhrUOvZ3wSTw3JbSo+eIlmB44yXWtlvX5zDR5UAD
Foxgw62uT/hneYIXAWPYeiiE1fJqIYduLLkI5Jb+SZaYVsAJrrVqHoHpEiNpxtEngwhKMbBY/lSl
yI1IhfxMV7fc8txo/ma/e0ZRK2m8Sjws1M0fPmaujDcl8GEk7o6ZXp/+WcVRTvC8ojghVfc/b5U6
sHw27P/O9Cj442vyZrzlVoWrfW/YYCDJolSyGMUTrsbs9+YBM7JuX84zYBl68W+Oq56TY5Sh/e2r
YLQK1TIFcqLoQZqAu6D9ZwmpiN+uNT6fNbPUvp2epNHq7O/JrQuEzzu+tfstLCUnT4yu8ZqUyuGT
FAznsD8VImc+F8eRbxJXLNyYy1bDwKNa6/AQUgpHWt/FXX7fPH8KnDFkbMDU56sZtuFx4ubCCAb7
xTKkOcer+TXQwf19e3z6h4vy2zT+hk2BlGGHTRAM/t755zCtXUYJNqWtJyLadsi47PwMVyDSqNDC
ck1zxxDOYNcH7Z3J8g3giTAPBNsww4y4jstZolZzOPTvoRuI6j2HsumSVgFXeeecG/SYyEZiTFKQ
22seI20fwI0Mnt9ISQ6ruDEyvGWDVe+Nd/1ovH/3/O/3bnWX7svwSF/AUzmL72GRMrVvCuMo1Ica
A2YXzYT6TQ91JI4S4o8ZMIcmk/YuJOZiVmFfSJ/z1FeZZKHuqs5wHBCAEzqCGCYFkEI7tWOiToPa
C8oElQHPaQYuVM150/dSvvsddgMhdPNkip7Wr23y4EqnivdY6wFOpstSaqJYIBdWjiEFSBSk960x
S7UWmC2PuiNJVHZYAaIvP0+7ElDjHulJAzaXR0Zn2J/oWDf1CMqBEu12Pp7Kpe11uY9iTAU8DklK
5m5EPB9zRvq203l04XuyZorY0LyjokKfr+M1gL+dzRUdhywRSDmfnpJGrLl8VpSl5ZYOM/2bQQUR
nO0m3UH79AxmciNhDY41QO6FSmr4GJV/7dcbK63R/viOPxUxEjqPgkzOhZD8iNoYDJVwYzxeQU3E
ZmUmGUj3rhvKsTU6i9ppT+xLhRL4Cwu0C/MbDgDI/cQdXLrYyO9FvTx217l9CD+AYHLEKotoVUDl
F0tSIvQ7z67YcU9cufZ3sTKTEtz77/PF8H+GIOAvGhmbLcFrAX/1zW+K/nJinV0UjrnG4bAAuVX3
TQBdmLY0MHzYR5yOb5IAqzcfakzroBRz6flo7WRr+sB1rO7cQEib6CMoe4mUVMB1/Vf7JKJs15E2
xllElwXEl/hSDrzEKJeMm433V4aQXDWuWWU7XjNc4rYw4alco5psoZXrGkIKGOErsoLzFxjwueHc
Z76yYz8e27EjwxgxMfq/tPkCfWOWymDrLE7/sQcAOXUmyPztfDyZ8NcedCF/5inYX1f4UyDEgVml
1Zhqb6rPScVMvd6lsnIu9iAjnbyS6BmgCfQzNdeO3+bLKvllgC+HttT/3SamZXeeX/NKacQ5ayEX
x39GOZ3ZT9iSP2Ig8ngDgD3CSXBtfELJR/DA7/Od9tSg0elwy0SEj/8apeMWsrLWC3NiRdILmLtl
Jp8R4u7BpvMBz4+RflHJr3E0nEu3RBeeVTcWjcGDd9qv30cDtNAB5zMIfORVS1OA3vOw56Dq02kO
XuuaybsAQPBPc8kNw9G/zHnOmPjz9Q4AicTNqK3kFT6I0BRgBsD0jtqq0OgWhXEUKwvWnhFbwHP3
1iBhDWb5LS38xiXJRmhB4A8X7mDSEO2uTaZhsicLCeFYw6whJnuuF4Ev/YsImPBFBQDvQ4DqMCbY
NQcULEQnGhwaldeRWqIVEOsxgN0G+7naTG/HULB8dRW1ikK3aNbtQI02KdgKNkkvYY/70qBx2daX
1+p5foP/TcDqu6nErni2DqENSF0vkx5CaGnYbLiQBrYyl/Tlpa4FVeDA0JvUzVm3x5jGhtPqBCBB
hXlqPiiKaWKzNda1waLSzOqvuW5CDzxeKZcyp60KA1KVEztbJn8cox0CDYASfTVq7gbXBywrzpQO
l0sgIzvxtOteYHBCaRhqo1E8Qlho2j1miWRnGG/AqSsmYrzrl62sLg7jvg0eTIAAyqdicJd7Hv+J
lROTbhVE+7socMpUXVZEEH6EM5Q+QdiZBmmJgbApMM2zj7EdYEhv3f38zsUHo9mlFewCln7dujAX
iVfapfqgSl/Pum69HWL7cikgaBFEK3OMZrfYUZSOuNsJo8uISo2iN/CiHjob+L+euDmPP/+4BUC+
80FFBhLgpauc9UMY+5QBImWKXDKp1dk6HdbqRWVxIN0s92QN88rSQuy2YZXgi6MAkKZUZyxxU5sX
ugHQXO97bknPHYCWYCSJq1UF1aZQiDuZ0gY5n20BoKx0v6xbxItO+dojdUFE9lU7IXvpf2O/IaNi
rj9Zjuid40FWcMU5pjcY5EOlvrbl33ipUHE/hV/SatN2SxPPE05trk5nE1sF9bidKEJdIqXU96tY
4Yyt2z5HAxpmfRU4+SVxeVEuqCMo+Kqgb8Fw+l10U4VoOs+nV89wc/WIlVGZjGyVoZw9hZyfAik6
/K/aMyKKEdwBJWoSNpJvd4KY+KddnGLDpBu434V13TxtSD5esHpdcY4So0mx8wyMn7r2daEDqQd3
9i/JuT3kEg/vAKI0dnZr2y4SWfqZKbHL6CN+C2Ztr2qpIg4sMbbcKEfzQe/k+KBWjRw65zgEnAu5
MtMTt6OaXoOLSWrhX/A/j2nRaGl3gBIET1KWtEjOHEZewLHp1DY58QR7rNY2VfF0ha5pYWzVVyrf
JqH/FJs1e9qgdEWESok8oL5lllgtWi/23SjZ0duIhJextiwRKHlG+RBtUgG3N2mriR8dCUza/iw9
FCzmOdbpcJ9cay7Rv2y4YNPL/arPZ+bYfe94LSU+vhLDwaqIuJ/GTZfo3eBncv3RNC7o5k6yAYSw
6C/T6VhSWvumjv8FaqdGalM2RoCj5cFEB0TabZmCfXbnUJQIBTmB9eSUwvqv2mKSv7VzHggIT5AS
I7+5I49/b3vDtyrn58eL6nbW0vSmH5J3oPlJX15Nz25w7XG3eJI80sTlTJAK1G5QzV0eZS50ckLB
ocfeatSv7giesaIbM15fUFlV1+lHNnSj9Ybx/OE69m3U9Pr4Q3Izacrd4JO7V/dlGgXQQB/ASbNF
6OopnQ0wE4dm5E+r+2s5q2Hs2cVTdy5jECbFzsgf1X0ZRnncDBaTS9vUsEbLkgPPTljYFFxUizKL
S1/j/csc5e0OfVDFJ//KLwDLuCKEFqlkKmFTGSdI9LDlHJfH3k+qk60JoBB8kJFx+IhMkj67Np+l
xKMkFa6f1A3tBn8O8YXWIizfN/yZ6W3U9LhTeUihMCld+EHT9SyQOjLn9DoCDGN9rzqCXtnGhWUO
GHKgslQ8gX2zcQWoJErpoMXLZYK4jQUEH5/9onmMfNASOlqKmxYCoef4EIkuc7E96AMvqGs0vE6E
kX4CNJYo+9ATr02FgRtDOo6DAZB4xUBS35LOBVHHi7HIUER1BKrUjh936jtL+oJTUj9gEcGZas+h
58kM7O6R7igHqXMVWm3JYxNw0fr0NuDqUsM71ejt6qlQDE3DM1Di2KJ7LRXee7q+3DRwJofP5g0U
XKtv3xOJ5euk32RLd/nzcmfJONVyIOMhJi3i4f9U5E08hi6dK5vdBrSHtkXAR1w7D+/ATheWak4/
gPbmC+H6QMNIeg85XMACLKseHp3r9CYjZQFlTA4fsOUx6JmEmq5pZSTxsmDC5ny/wtkPhbx7/f6b
S1dw+pASW4IBY5XuaKAv3jbfmGlykNbgwbXn18zWRZxsPDu25GGR+GeT3g9iNi4DaqPJxpbUFBex
Xs4tnOmvDSqltbWTyzi/TDi/T3ZaIrX4AYmi90T93l2HSF9s23h9aA/lOOsFdJ89l6GChJLsGZgR
XagkaU9K/vEBkHbI7dia9JG20rDdLGi6JvbcAeH34GjZF2o30OK+WspzKlugoeHOAxRWoEfrArR8
PU1FZZIS73nQFvcY2Cx4SSRzrFAkpCUGX1dOoOZ8v77JXjM5yvw2Lv4e3j/nHl/l/8vyvhXqameM
LPIxp09RtHlu+hCRIdm4ljfim8qgiyz/1CZP2zAZmNTfPq2gHqBoRn47T6651Eaae+njheXXtR6k
+1949ClRpMsHarq/wWYmgif3uWa74ZtBa5O9onifB5YQtla3U+KesO3vpnXXxNTiaV8t4CG8RGYO
xt0yAJ18uY1i2k87tYxyoKBiqJbpWRUGivNigpGU2R2Q9/lFCSulzE28TUwu2s3ZkhEmA1ronzKG
cQMnWRQRScLgVG4HbD37FRVv+384AFm82bX51dp/zN93+YKPcGseLpV6vDxsHInMmC84KVpC/8Dc
I/EHTSo5dM2RvB3uYGH2Di7L+yL1CqMVcRn86asspX/ADwsH8rNRt0WSzSkx5A0BjxbsjPSNRqs4
xILs1lmrVbzOpXYvamQoTADUGxVRXg7PPalRhzXtqdcQ6J4ObIFF6xTpLZYm/QKim3AInq9caSIB
IvKsSCiLF72y1YBJHayiG94RoPufeuafyxFEn7Fzj/wrk12J4VuPHnT94eQxQ6nEqNo0AU6Z+Vy7
YblaegPLdadhbrmE0KH0v96YryyhARb+Um63Pm1w/ZytiKq/7V+WE78xVMJLJ2gb1KwOzd/fueoR
It/xv+Dkft/iWn8TNHuET5Dv/aAGUbLQjFbDW89Ei3YtUgHLoILoZ7Z3wJYBnAhmv5Egl3JXybwg
ue/vld2qbZcwSputKdRg+ZWzxj+mW//jDOWmOHgWjWFpS2zTbtjyi73GmhIELnG2+x1U0ZVCoJwN
H8euEz0ctr+MI4BLQ1TY0r6HOot0JOkCBBp9kmSorwZncvoQpzI5tNRRQ+qx/q820OyceCT6qbYj
WfrSCsEx18wUBuUZRq9DefHm1lkswR7wxN4pD1qK3m5kDYPuFvCJh2SK4V5SNPv4bNWVrKG+7k4W
ecrTBsdUdunL0+GKyfv09NrQyGMa8klftNYi9vg2t+VBc87pXwnfNkRxJ3vgCPy8+8av10Bn6iq6
e369B2K1uHhhuQtlUWpyaaxyUseiUOCsbXtar70oYl05HfAB7ONOe5Yx0mQyPQWZgM+UAfKH6YuE
d/e79vqX4nHmhrFUVaKvORjosKBDnh0kTXRU65ZHoxVZ6NjeF/xV5i+tBP1zlQBQgSZkSZlAsICr
KPLm9lJzgJBqkqG1vjaqAaJOTthgoIUn+mCBMuV/ue5coQpaXDbg1/Z7jjtHYW/BweRryYQzIf93
DIl4GFguoMhWFlLmelWINaklOA4G7HQZU+GrD0hmCaKIgVL0QIxtKMbScXRI/2jg6nEgeD0N8FoG
zFmaowMsTjOpGEV5wi7yF3CMH44+1Qtck+uGjnSx8Dkblmdg7l3wWFJ25eVRKSjRg43pf5HgdbqS
NZyP2utExY6a7VK9GsyU+2R4DKZ3LDuucy49WJpQwdiYVGwLHRSlsBlcSLq8NHykxJKol45B+9Vn
s4qdyzOZ7zwTNljpHkwCo4iJXjeGwa1UUE+8uq6JGfQ3SDzXf5JI5HT81GktEYgcRTbPr7p7wv9t
9RqYkRhdpOi31giHA6FIN5jdKBys02WXigXO/R2irZQPyu700/HXn8cKNS0FduvXqGbDOHfuleNN
ieio8PmIa9DDxP0fAmbEfhHzyyNXMAA9bjp4zc27flnLSADggY1Q3Tz4zzbglX1VvhV85KByP/Fd
vZWMqGUL8DmcQOEnPbocSeYAGzEt8YCO92+mY5Cp6BtY1dW6mRB+CeOwXusZWTN9Y3TLk7UNjc2V
E59Nt9D6XtA0IuD7T37Ty50rEVtxYK5lMSX/QD4cpiT8pdVWk9Nk25mOd6pslwHj+hhVHe0fbIXE
/tRYvmcLcWWo2Ose3m2YI+q7g/qCr2RsYkmmXbUBDTo/T/uxvRevWIaXZhRXtSG3LaxsLZFbenPx
DiXtsii/KOkng8MgABL+ASHC8caUvw7CPWdS9Qbz/IG1y5CMxbibl2QIOKx03gFiLemHr6oGVIUx
3gSs39fnitlxSyRGPT4iT7midBmjdoKUa7Vwjs6Ev3YK2nS2IWu9DG3apmeSkauuhPF0CP07+fh8
j7ddEOI21Y7kc2ySPuW2BgqhZZ9+o9uj1Oj7WteH0VRhGkCHmAOMLLQEFeQnvSClax6+1g93mejs
Kqgum0vKLS1UGUaxfwSAQBp3ih0A4OGF0Uww4ylhVlj9u+B0HF/DXbuOXH9VbReExA83cVcg5/4g
VVBjVu46EZCFQHjTfW9quXbWnonUMYbJasTTArWxf8j7orNYnUmjfoZhXTFgCyBHISrsvuhOnR+Q
ZYHR29fDTo6kcJYHN5/GY4Mw/dqrAjuZyWpX1rPLJOPNqrGFKQkLgamhN2sA+yiX7XPaf8ltcoJs
sqncvYNH6lBpYMF5iswcY40FsGdS1F/faOazoM86+9xtCvZEbG8DNKVIeTevH+VQwDH3/voazbPb
qhZJXmEEhNCeAtM90oDuQUd9V1w3OvX9exDLcSYsroxmT9WkWA0Ggrw0pSRtGkrdegInFtIMATzk
8pvwViXp2acRpcRgdzSD+NkTJ0nefEQfM4Ub4NfkzHju4UyQAP15FtOH9cPmjKziiE+Wr5G3fhV1
s30qBUHCUyNCLzdRGW9LQa4Xg5J9wPr4Sci9OtA9iqZwS7+8HfGGR6yscCMNYQvP5L/dTssEVmzI
jSwnD563ly0wo5xaP0HGTDljDKxI9GGVq7bJzyjgRr6TXzckSgOHioIEov5DBMC20z4J6rbtu+lm
0Ns4AljHk/bzXgIHLsLDyBivk4yqpk467obrR3GZy7EGFMX577LWWQF91sASoieKMcLE2IdH8B7t
CUWf9qQFzSmp875opRSomEdt+o1/tstgI3GjqDOpnLkCKvwzt+m+HU4H8RFJPwW9iAD018qkFfz0
g9opTSn3UwU13shLbZtWgxG9jKd+5ffK+YbuVd3qujKO14RGvPavn5iGT4V+Vgz5wDTwTnxUJ4y7
wrKDladpCCSDphUlGyx+FGCSdXQ9OoVYMwYPOTdMyu9KYQaXVOyHQB1+aUjuJfepGnVAZNhopdwm
zOEvKMjofHjJ38GCEEtRREGkoRttGiZKII/e5HFqwNs4Q/7R+tkzTsYaKvDNCzEY0vgq5EWFXCb9
R/BZvBeiYG9xUtHBp0YdUlFGRf9DfIKSyX0Oje6b1cty1vcPdumxH0t3w37LSTihEdjXSALoqE9c
7+RXATWbdoXBdhSyt3iE9HwFXp6zerNyxDq8cuW0GFovjhpdxxToYvPR/86Py2WubpVMtzwO7eiY
ksYxSxYm3QYeAycmLWiKmGRV6QOs+/dMDacaS4J2pq1vU489npOCe9e9WbxWwS0dBid91X2P4OK+
NfSaLQqyWufw+sCp04uwqyInaBXdMAcCl+BQFIfK3yO2l5vzmCizWMR9zRMryb2FN/XoSH3s3Pm+
6AzM47JarpV/NXDkf8z/wjDlB+nNO1NGJBwAT0fpv/Gn0bOqC88G+zrNVX9MmN3fy3G/I29pmZER
uzJaShsNpELhnEQYOs/w2bjdDwlEOQq/gZ6YiIbjZmcBIpXwsG36mm0BcJEqG3lij4+Z6dkvckGn
kBoBrbhX4u/z5W8ItGx4GNUakHtHkQuP9cCYFCa6PxqlJ4SXa1LmwUMasQmQxeWL5h57aa3N0ezj
zc0X3xq+4zuzG83w+90KEeWcGmBn3sfvMFUpL5iYqHv4760omoCJYRV1B18KDArkjWWcXZgO81GN
e7iuvHfCZELdGOUJAd0z10C/Uv63mIWth5xcGbJe7WwIoCoMCBP8jz8ZtG5q/aI4R2QvTKV96Q6u
COKgGTECwEPmO2PBtPh/60Kbe3R17zu3+WX1NajOZtOMjovwQ6+hxlmZPj0j3cQWbvZaVbwf3Y6O
ZBRT7I9ApxMGcXmCm2DU03JUvb5AUoPoXuvy0jitJcFakHeOMlJsF0UYOHskkXW+claDiXQldeF+
O7LSH0flV6pzgZQMIEJArR2JjNCXcN6BHX442KtQAn6fXEsjrgifsJV4wRepxW2VfkxCQVHNbhzH
2DFIQMWErhx08xCFYsqVUK3qEmdx7udFVsSE0p/egjAx0oPw+PdgFbQzdGPWFYDdJtUdO8LcbYrG
jXmrelpr6wK+T2muGJuril5lP3kLQOb7tiHX91YrercdKysQiGzQPr2hkzlgONY5yEhHB/lpDUk/
b+k6FLNBljwWrqSuTvn7hCeIDOQ1eZnB4tsKOGFQETAKmh1zwI+HIduHziSWIMLH796vdaJjd11e
BM1qJbPtS/SU92bB3AAjtYKI/NmmxsXLyxywXjdYbemVtM9qpHOtEpbJtlbURfRBTpNc8RA6Tsis
aH1OlCnnu58T8pmPH1qsHux+vcXWOSZ5Ra5B7w44Ta/50snyrWhvglAJDpWDfTJrIkhYOosFTs+i
QFl3umnTfFXJn5VjERPCxCKH5FO4wJzSqdmdMSGEFQGY5Mm+Jt/a9TsC+DisA6Y9tjnaqNv7B6cj
ho96eqieQRIv9A8A+t20YjS5jSyVCatkHDVR+Wfr1m5AJaI/V0Yd+udJFeM53YfincjBiRmUydJb
66EMrHUDnw/LY/COTgpFTUYA/qnVtPG0p0kHpVnqgpJNzNevZRN+SpTpew6RvqamayAF7XKhUe/c
/X0XP1IMe9u5cIbvKRow8mwp1qhIT6vElHHQDJJkwpOqmUYAv00Ap+V4CPWazDa9i5UgYH1d7hRF
0MlzPDttyqGGg3BIywUjl8sZ7MPCHsHJefoNHkS1h50j90U0AZBC11eGv1+yMKFJnKaaOLCo3LoH
MCm0SZXN4ajfaYGGge7kIuXaInvh5EsOpKxfWQjF+YEWyLUTaYnIBsuR08GDbXENgEyw1NvoELVH
AIKJkZfgti1E83ft7Ycr4rCuHIoBtuQY2vcr7EiLik/d9p7R8+iNdRTeE9JyEK891rkdG4G5vjIs
Wz++OiXoJi3XMRPnAlt+X8FnHxGSzOAPDCztxkLUjveD7H0EQINX6qYmDVzH3S8KlLpEz/Oak+v7
U7QGBZXnbNj4j7uSGvl5LhHpPwjNDN51njMwzF3gzD6jbvdBpIIU/6d5Uta0difJVab5BD2s4FcQ
hyY68RVZ1Sv8kqlfhbn3XfiQo86f2pA/jwH/mhboJF9x1g/bxJr61cGS02SdFCN5S6avXxkATxgA
7836f85j1FRlaws6dmUbi/YEiWDel6r+B6TYjQHdeJzvKUSJKPYU2YT8lseIYwah321m1tkrzcgw
S1Ds4ge86ifnbNhLMKdKllAHgyDZFNqlSaNr614Mi1jy6PcUfpYaQHomTdeXXfI9Jzlze0CxT1MO
cDMdSlYx5liKlzf+ujb9ggb1ytsT1I4BV+6aMlaDq9/qy3zXvYJMsWzGef2Pzs/mOG0E/kvzaQla
Yaffb8NbraGeQqJ/mcUneUzFCBf8Pcmt4yZWeE5bBsi78Qseny/GWlQ+IKC+vFSbsLx9nzfaudRf
sbUG0hG5MKoAu0+qtxtOvZBwKi6ovu9sR0Cjb0+MRDM7NG96zYIRFtiswGn0xuU1bNsPuIVr4SS8
zX5EzdvHu7Wt5yBK3wACXmG9CtixRywKUBjQwZQbCP5tbBffQ0Pv0I0foImxs1MfzdUqELOw9RXt
2Dng+uRS7AOdkXWlJBVqSN13AKn4ibxnu2gMQNZGIbC+OWbwMtEjyq9oCRQi3BisfRO+VfjX1/JO
tusb63RJiq9Xq2MelhUNXpOCrXDPiNGGkN69WS13/dnawRhsOc1EQD4mbmeOZp0roPbJY6Qlcphv
nZvDJ05R6HikRax/7NTh6kWh99Iy4pZwa2e0AhPWK5UA+y637gZvFnMrBcwgozGQXnDP5PQemCdT
oJbZyCB7eSFSBXvnfBYA4OZGgPCZIXwGt0ovUeQHQPIdQ9DZt+FaemcbaGfbai29I+rh1tHdW4Ib
CplJKuj9aCt8eb7a81E0W6Q6tuucw6PnkGFMty16ZuqATlp84HKpklzsRFL9W0/xQU2pB2DQ4NZm
Glsu51QaoTQlCNbYLIwuzn7dQzo9dpIzO0KFyaON75Nn/jxMR5Fr4fPQa6bvZ/PrlFZ407wKhdJ6
qjLBGzqXg/94KiTFeGVhdGSGTOcI9hBx5OgsZ8hQg04VTCWO94GouLQcEJ/vTkwTrDKU5T1SPgA4
RhQJ4H1D6emYf/y17Ld7TCWrA0QNDRojha1eCNYWTDJooDvO8kALRN+yFwoehjgfrlgNBpzJtEVY
e2+rn/cPi64XR4uExW66eav0TrMaG0Ftvb6TSM7SXMcffnQ7t0J5ojxVihMUAOIVyg9T8eiE1ZqE
WEeGm5QVwlDCSCB/y6/jUCNWa8rG0mNfeAJfb6A48V3DVYYvpjVb2ldJrkTz7ZplgDfSdFxVswTY
UeThoAES2CFTIlMAWIhUV8RkRp5HLkXai4FbFOxhJ/XfkJdhkmZLvG6nvanPzm3ccZAsI33dxmI1
Hn+YjHue8VyERZrhTnHnba1US50LhhqQx7YZuujCapygvgxX8acwf6+pbgx9ZX15nzh0mxUJzDdI
BMIMEeS/943xC7jOPYs7u0PAbn7B+9HnOcfleaFkvTaqTR8yGInrsjT4xxtqGueFlOXZbQitEEnr
WRE8cuiq7DhI8Ae9LdTvh2AE6tUurKRBB9Yc64nvcf6ZiVmv/YE95pN6U6i4Hg4KmnmMn0AjRSFA
F5bNYWCv69uRHWjB7ZI4+aWQnZUKuwFahBKQsd0Y7AluP9/dzv/RRwypKmwjD7k109zACBkImmXc
Xk/APG7OCEqzVmEkCFbZcVwYDlyGtAFZf3okDqc5BqotxvZ+0K7lGXZ19aFRieyaOvxv/lh1JIT/
8C/dNQOA8pTHmtQw2GwNHGb3//cHRYJRDG2E56rWyXde8S4QhnWiUFfh6NDACL0TYelYRjjbpKsv
y/c8txzv3U/XDSvMzpjh4KjDiG3RNA0UxknOAW7DtPfrcluEoog8z+DGdwD6Ucwh2G1CeJ6m7qiK
11rBMjYpQX7PtOX/YRANHlDQz3/Fy9SJXebk+nnyo/lirO9gux16cWUMfO6z90OYjK9q6fI4XZqq
UefU7QPn6sT8v1gc8E9c0wDwJtVFoTPHOC53kx25GGCAkGmitjxLOAQuU4UXlFh1HB1ntOvXzDmQ
erf/wb0uuSt5NJr6oTNIlmyHexT27hqVvOYoGOHg9rDmMpkUlqzPGUhLjwrvKoD48am1JDwaEdf6
9N1gy9zE2wXc/4X48Gh6PYVh0fRoBhJSOtsN7L81JAoOjGtAUwj9NV2hbnX2/SqF5K6nGEaEq6uN
rvhtySoEXijr9kUaP9/7mgRarNV6nTWZkdO8B4YyXAdvS2DKw/43G12bMKOn/h0YRQGd5Ad4fl34
099OfibBnUUsSi4VTfpLII42sktO2aUvloWyP3Lhk45lpm1eq107SLDyFCurQQc6OGvhJggHnG48
I+muKADUWkfdhQxmOUf6gtiRUV5Dboha122WmBTX97WKnhejbmF/IUjm+7vNfTU0EygCSBgLHNAO
q46I2IIPlPIWbXTwKdomB8/gNK/vj5n9wkEYKTZQc6kavMhugP6bu5CX93yhtSFyH1xO4bIkgr4e
pbQlO+Tuudqo+t0gfZI5fHNSGMcvdJsBgAvVRm1wZPCuTg1OIV/X0oFsV/KWYDahzX4R45gbWN6z
AXW0eq8EjCxKlxKNPENP8jvTRhAHlxHHFWq6defl1WXvTKlevnQXPd9hymFrZTtSUYRvSex2cX0a
8NSnvy7i8kJfNFQRFaBRd+ComASQVnMC9LeqtpMQk71jxrGKCsrFM8lbzhyUcBj2dkTdJCJe0cSY
/LFEP36lW81lO0DorjiNR3QdBcgGBtwCisKCo5bK7iWy8iL6JA0i/FC//BIn0YrmEyV+uNAg1aN/
GEhqeFjQ55iUVrs7zuNIdqEZkyBAejdzRc5YwFAG0NW7aFWWnFTbXco0BMNZZzqQ1kFWbPWf+Imj
PmKrDeXdsBYn4OLSjJYrnkl5Q1UXBkb8iRHuyH0ZaRHGCz9RDJRP6YVSp8ZmCI6kWLukLhrmYD1W
MdRWLHMGltyIEMtK22mnrTsr37poE8HB3zQ7yhDAGvOmkpEuzWPhHPZ93wnFVOLEAPu/qrCAnj39
ETR62gh+PPso0uvIh0XDApnZ6DRI0crtFmLPYdrQYIyVzlW38bAyE6T4upjQF9LtHl9qjD+KYhRa
T8isugFFGceG1JEkHcI3PRoqgSVmI86MjxFiDu0TNXdGzCh4xfUkH2JOD4NTlXwDe7QyUsjw2iPQ
Odja4WU7t36of0eGyez5PJBNJ7AF9znjYJ44mwBHRPoXJrdrjK8IuzG05EA83N1s7dTPs7s7GI5x
z85vC3HC/CE14jL+z/IVJxq+qQ5LkH1MYqpUtUd2WX9ngpIex0rM22+ciNdPn/mUztIlJMrh6n40
4HyZIxsJV/BpCeSKxJ8YZnuoHNBKDge5ZO7p5G+FQtO8QTGg0R9KA/EBsZ0mOO82MkMLxRvVU77U
QGvN9GtAdbTYh/gpCjviiRAH6Bgci+3Dk+vrtL8wXVEDAEcVGqNyKABVwvKER0pe1zfCUl5MC+MR
Q2+3yIwLw6/Wwkw8/eWXt9awmuw/4WRV9Q7QhAefWmim5Jv9Puk8E4yq+TJ+4+VwTNBgBrtI0n5c
IIu9xIIn91dkewz9oYtHQ2vko2LS5tI0EWNW0nBjjHmnlpSF65Q5TjHv9rjZasMMs5JnbyQLasXj
AJV+JQzOgkCowwVjbZJJmwPt9a9o97rr0HxXKDmQGRrLelGiojkamakPZdG22s4Vb+D2bYHECpxn
Z1yH9IHIKTLhOlVKrhYqWLyJ2tjxe0GxydikL4TloAAKHbVwrghJxpDn3sxonhbMGoPNNOdeedrR
BbrnUlQxID9qXao0NiEzlZLqIDErtx8ZS8IkNPKZWhorCb77peBDejgOgZCLNzyknjGzFCWcamsp
YLItalf8l7mcPU/NlA0XLwtM3dckz63s2nbcYu7qLqaKy+minnM3IJ41KqUJL+FzhBs9jD32wQye
/Q0atrWVrCPZjDbXOzW46NbwMpaBKq7Zo9H85/ghYgTDY0hVdxZpPs6Cfn/Awz8UrQItegqMwwP0
I8IPg+bHVK2IlXZK+iEPI4Hct5zy2oLbCDT1HnbxZoa1a3yj11AeDVtCgrde5FKkGBm75Ew4ugDJ
WFhzVApC9WKXzDJ+Ss8Ai5/0MWofY9p44ygbe9TWcsrAMWy1etex66FxsocZ+OwWH/GSP6S6yHOD
ar5sCQDTU+bQVxhfU9d3hVWZJ9KxzMNzDumiVJAOUVW6ozJ5vrhdWjimfla9dWGSbDXxh6INzGQ7
cFaOqowPf86ocR+3Myizwb1tJhHk2lv/g61UG3pP2ZFTmwddRkq6foTvK2E4WWLA72Baozov/N2G
YW1j4+DEIya6Fpt3C85ubTGJmaKWX+nJ00TYvSF/x6UC562l9atCTngUkFf68YUXsf9LngvA1t4x
1rRkKnXvdjM2VbAnA54mXjB8/TJL+P+PVx5xEaDAKyhEH8uUAqjk0HxWfyswgdzVHQyywASGbSWo
PhkxOZPnsCJYvTkYhQlJT0lQGafgy9+dj6t7vUxrN3cqu0/WCbo1M1+1367Ve6WHcnw6agGFlpdk
l5OYO/4UeJx+i9aqAbuzYb+F5sZUp5tMNvoLLR6Szz62Hcasah0zpCrEXqZhKjIqZ2tzL7st0QHU
xdc5hSBs4+eMDOKTRd/5J/eju/G5uL4i8skCNKd/O3xJKN3SyMYk9Ehp7+fdRDwcFrUOM1IMLyGi
KMUQwJvNlUtNad6+eDfp/QLoi16G1tmMxdxaF2I/9YPsOqPwcAHjCJuiUvz3LNoWRR9whFZjEO1q
sQCGeYDFDsDlSaXHA7e3rwODpEIBi80pHt10L3h00rrHc7oaOhRufYdbOvrCF9oZygfylC86F9d4
FydeuaC2DiVCUslMhZGZph29SsCk6oZSLsKp7/KnIvwpc9DAVeAiEQ5J4KsQiQrBZ5R+xXolasaW
e9m732qjTWcP2EbEMq6XdDuzHJL0QtL15moswU92ePoC+Vv4IouO1CYP3d9+huvezSjg+fBeXRnh
6Rx5Pk1aEGhyR5LD4Dut/eRSA/leZP0XILQ3XEjX7LJchOW8OjhcIZ/LoejXVvJ6KhoRssfzPkaw
BmvtVowWTgzF5peUWwFpK3bWbT2CMIiUywfJxakPNbHaas5hEfB62dgJ0wF0Kh0dawdYnzRSjzrr
h5/Iw9lq72neefw18fOrpV4IEjozltTV+zW1EH08ilblFmOXew4ssHtsFd8V3DNVSdTfeujgt1Hu
HSwr+HJscxYPW89V48jY0HrOqs8QMz4JY9aOJW1wlUgn5arTVPehSx8NRMt7ndPZ9adWF9g0utS/
nZ+CwMw7+XRD3prb5MXNPTQfcvBLWG5+pIkfzo7OD5nUVUon8Snl42LdHzF03Y0wANgp0hOb4dq2
qxmotRmtItFjGmEG9BG1v5agf2gdzghY/XEh+TV+dyk5Io49nuhtZlzCnY45MTJsoh7TaHMdXf8B
JkXgOLZYCzpfP0Az+OT3P1Ka6JGbHli+4Su7KmumvlTy7iKA1Oktfu9xnZkmbvb97PIfe7J+OJnC
lF+M9qzNk00/h9ZOP0nSawoGyfhjmT2Rq2MRzVMj11usBL5kON6bbzwSK6osNRwySqYeXUEWNS4w
I7Y9Xu0eG4P6GUr8wpS+UmWHp7j/Ith6gGN6oyXeS+bYilV0GRVPRUAAT4uuymByJQSd6EpEmJfn
foeNqQna5wwbBHqplb+PFwPurNWinh3T6daOY7l/E2D8Zn1duUhjAYghqGRYlEVfQjCqT4YgtL2L
DbtfDxOd3bKY0jjBqAJwl/GEvDjk4d8jD5kVyqBD43D2fhDIni9Z+AYvcACFJs5rBeERbTBNTO7e
6VEoN2lk2jVI3g7HSfZT2FZnoB9iQrXHZRqrN/DaafXRGRR+ONeSwVg8F6+PmMN1LqAPS7Y/w0+d
/eD9YKRvRySd9Qcu8sbG2tYYFyGsDpV8VeGGCi3Md2E6uSs6ZRp+GKIvLiAf5dDqnBdGPMfQCDEx
rbu6c75PXgSLaIUdmnzj+hWOoYMfHxzF6pHQHZJ1tevjO+xCE9p8hoLoioNx3KjEcYkYClos+SpU
WxNgoLOw30nosceU2daixgajI1iLAOTg2n2i/tzdSb6mJeD8ty2/Q4OHTdh3t0LcI2wfkfrCX+1Z
P0/dd47DNiOSRNVfN550/w/21BfRAadTSMjy92b9yTdq1CIBjFJ2A4bZMG4/gyt++QlmJ6iqS9j4
ZLNbG/EvkznByemUZMa/Znt9occNpsPOch+aSnVI1moo7Rp9jYWAijzskeKHPKTAdDiaPxW+NrJX
L5Ki/CawOP7IsCENxbiCOGx6jYUMfJ86xj49aSon2phagBFA7o2Ib80Bzv0SQxTJOBT6+5bJTuXh
8F+CZZninUmKPn8ZsUDn7JdLtJRulQ/WoKy5P+U2DyJcZcCJHXS2BXGAsd33EQlB1ZcDS3HZYSN6
U2NZ5TjVrdgZFuDS88X/KINgKg56Qx+jj7AeVx3LKKKjuFan+u6jbOL67Tl7+HgBSQ6E67wwIXfb
3MqFuHt8Iw+VD6FaaNcfw9PyJKevdSNPYaBQmcYBr/H7F1Qha4Rpk5Z7M9fgt5usjs1ULbhF1sVR
xkFnvwadNWhUoBDQruV69QI7o4Z2SG0uheIfyVsmaxSW2PrcE/0oTHd1weRo86xEN4PGA/ly19fE
AOjP+w5fK3vcaKdKJGAhfSPPS/kvjfpLmuNwl+h9EsRWt1MsYZ2Hj97G7rjE0KFQ5oHXhW8TdweA
kmJHDLmlg815RkuNQ5xFPM0e9DCq9OeGdM7LFiyj185KYFSlTSXbPmHt9h30DDdfMcVIvso7d6b1
8jk1DTYDIRbYH+b8FtMAe1VdWxNBXPQvHQVVBzkE19dDOXoB+eEh9uSYhiwFFRkVxcqEpA/dPRpk
cSprSyG7dwSx/toQvyAIkMfGfOVg2eBzT+VJz6oeIyQUfiUFGMOrT1tBvq8EhNepib2UoU9dlzEr
mp56TcMVewd/Gpo1USBdvttGw7rTZmJtA35r5tpENCF+I0lZaqOP1KhV85ZIy8SXwo3M7VLegtDN
QhAXylTkJHwDwOMA+NyWp+kC89uPkFEO6YqtMFDz6QSKBSfoZ3XlFd1JUoE/hvLdbY7P6Qi7UMWh
XfK3i6hQol4xnNiFySf581B1qk0zsjn2LLWLISXl4xMsREnURc8H7lhbR8lM93r+C6flrw1e7kaW
xMIZSscgk/n0p/dgigv92aeIcS+SxS6L70dQ/e4rTHjkNm6WhUI9yj8JhiksBi4dJcfYqbq8uA9z
v3AsyavjS73TquMCVwSyxldFrokkpqX4WEMSML4JF+WWN2T5k1grQcHQy+CzPkps+aK1+a1l3JaR
MAM2BiUlRMbHOAkGz9GBmYiTLxDwjk6bG+W8kd/2zoL+lRZ0DHpwDRHKsqx5kZcPrRcFxpWiSGFB
6HW2wX2vQ4n60v6dJnJLRssZcknHf30jfWjv0UH66letpP3hBOudaXYOgDFVxtFC1drA5ayxOQlH
M2nVa8hEk+/ermadDaDOPlxI5oliuUCfsCKtO/lE9+nSAxxkDplEg87McWo1wL5P4bW+8we8RW72
1jJnejkSqsWB/kYnctsGVXzZ/GsyJ3hwjtAqWmE1cZdzsGNBO720JrnhhXkQli15Lpr7OKo5a8wD
Bkf+M8PyuYePN72K8EsRse7o3tOimQ31CsX2fGpm/9zGpsnbqLU37tCtSBI0Mvu9mgjaFFiN37BY
zF7fw0Sw66qxcierbs2dZ4uWqY2Z4m7UZuebnFLF+tC8nPyV6w8Mh5uAcsc2j2YMOZ39CDnUd+5k
ga8KIq4PYVM2Z5Q3KaOOCFFxZddNPINkJwk0GEIWMhBC3SbZgjF+EAHf1DflTqszch7UIJnKpWkJ
h9CjXZaU1VviTjvVwrkXYKKsi6b23RXrxJ2E7gZoHfRDCQqEcdYg0+qO2f2BscahD4BMygSnsCac
SzMoQnwRDKOZ4mOuGt5dVZ/sEbQzkI7L02qBM/UYkVgwfe3VAVbkTaaUblt97fjQrMa4/tvI7DFP
JCon1Ks/dx/YogOEQRv/LCoMUZkQUKFWG8+C7AiE418WdptJB1C5bxZJj5fj7sPeknBZipEU3b+i
hx6EIhfnYJTQsA8KB4KlBLCcsPhFPk3cpAxmmjIadYpfcRjk+FwLEJhg1G+AXYISuo/Mm+OyCpXG
YIHKUdV/Eeu3WHew9wzxSHU5zReyGAzUiSdwUVNABYU8VwZ0nya60G10fwAFECb5l015warct+dr
7+ShmLuyjJJkSoNDtkZwns9DTS8v/yKDuWDrwnD8hZByh63iB8MlJ4udCOeHW2xvvjbwnI+Ahb3c
auSNg5rR1Mb0qpKH8aDHecmd2xIMNxnMDHnE3EkZi/e9niF+BEvS9pXpuqgthSDH3b3HQBNAXHa6
DJEraZYCOLCQHAU0VHcyKnREQq+NgYcEcbb7MpFZoJCyRPftRBZalsKcQn2harE4vQUv9ib7gI0S
3XZDXWLSFbo+pBYiLu66xrttOgchCVf00iXsA+a1J87WrwkB5BuuZ4CoPYYuT6DFJxSZkvMJ0QLM
zOaDi+z5mSGUFqikLbmXfSnzFHJiopEmNpq0CB9yuZc5Nx09Y6GyVOhH40l2q0ZBrFBGAB9X+vjb
mxzoNMcWogcVlT8Ijx3UsxzTMZ/ckkzTrk9V+vcjeNt2jnjgertYy5okz2c91k6OqMT5Lkm7Fry4
u023+9tMTWteyhWk8T8jcdv091XzsoyZrc1u8w+5vJK+XHXfZkv+3HL4S+y0j6UGQgFqVqlFhZP+
U1nE6N9ou4ryo5HkjYdJwKXvhq8xvwm8PGpURG8l3xjy2c3PLZXRRNrmF+3cgJMBhd7oiY0e+aKW
Gz986gKTjKHmoRWV9516Mm4AfGWB1ZVrltOC7KvkqzB68s/pw7JpGZLd+YKqyVqwjxF78LGVfIgG
HBaMT/J1+IdjiEnXognMO1v6lRNXodOlgiMIXleF2jy3eJu27yARVTOvdiJYVZna9mSVXzvdSCan
UjTfKxDK1DrdeUGj6L/95NyYJ5On8+Xb3xrlCdHp9tUlDGb2HjPpyytow7pvxryRlZKdJdebaJFr
E82l4AiWZNohr9zi8k2B4moA3NLraF8RSc50g8zseVt+FLCSgdRDRVw9ZjEpevShpfSTjHnfh+eu
SJorVKJBTMq8TEKAWQM+Klpjv7Q7eBMnachn6pgoMugg9Tc4NMFNEOjLlLVCsX3rDRgfyeJDl4yH
k1k+9+nAsxV6qn9q3q1v/UEtf+JuUKLkbpy74Xyr0T+d/tn5qtDtL/GlqzcGs9PBHCvQmWTTBFzK
ljWGJRn22KTFQK0X0A+dMVbdCKL1CXoCeQCylqnLUyR9yWMaOPV46RRDxuSM6TY0YVpb1k2w/5/L
pYoe17ZF8yLiU+IOzDpYxPNiSeXsTo+ctW8MFMhL/OVUw1VMM6gCG4paLiQ0yKvFf+vzDV2ZgH2Y
vB1DXI8/lCPoy38bVX6FHBlyz2Qdn0abOLO7cvXqvEU6QSq+9X4VyWEZRVIFORAZvzpxvI99jf5k
OpBzkRZDpLNbvvf0UuLLjMPo0a4pPXTjdU/G/7HTZU5hkXjQqPw9d6TeG8ifzP0dI+DFeJCh1CFD
yd5Kem3Ooj1ZZ1h/vcVSXC8Pnb+Bt5Nm8/QPNOfkKdC+z0iI7UXO8Wf2pcqsy68dKmTfmTHA3ILt
fEV7aElUNRAycwuVK3nlm+M6DHxohavZ/cxWGD58Tlv257EZuWSJ3/8e09mbZCHOn0BEcPqccC7j
e8prPPbBOBLUU8z1huDGn+/X3Ay7xtxpC4OCuJxwKXYvtU3lKdsOY/qji5EWLyFsXC/hTBOsXWJY
SQRFksxGURgy/At8SEUvgCz+OOZXldPgkV9HXVZ0BR9VYxj6KwFlVDplAnC2NMU1/E27TnmwzRYy
ddcwZl3AKFkVb9ayCr1YQd8Wcges+MyfpodxkzHTEi3EsE4yznHmYMnBn21HzcUDSfXN+69j3W7+
nwfkWgpHKZKzNqWUiU1KU7u1ZC1Vkvyr1W7977CfuQuVfv9GrfIP0llC7N+ey2f+QWynNyT0Of7G
xRcY0n8IicooUDT36JYV2OJdTvfep9q84avJSFHK443gAZZu+OYDIQk2XfiaY90pRcYlTJk9u/5Y
ephxXmEsTHSF1xTr6ls9KgqULzVj0Sl00/Xttpq4+rXnNi8S59ybsKo+rMmG4PubJjZ824ut7PLo
4KTOr+uf8y/L8wJgKMyTpdsMcw+wThYwECoTe449SxV21nengIvwCCtVVS7JmnLeUjutxzv9zTYQ
KVpPFvuuO7cgVcnUCyoyuJbsNxTLJ5SkhNONVgca1F08UOhoAg9xwAAFGhBoxJWzyepavLi4w///
g4FetJYGtvNWprQP9js1JYu1Kdb6wSrFRcBgzyCu+TyQj2a/vUWCcI+wCvYOxTPSEquAKB7dNn4x
s+Yf8OziZNCgvdtQ0ncYrimiKvZNch6p3m8pAO8iEAQ7XXgNnDsOiA4XkC1B0lmt3nCIG2wWFHp+
TyJ2mtSISbkUH2Z+CsUdpkK84nIQlU9memwRKyS2zDJHe+ho4dgtLUXiCUl/29egjSjLCHbbMUo0
j3GsNbpTEPHEX6ox5DUdfJfwsKR4DJLQjQP5mr7C4QcuNg0x6vqM3Ny+oVWsPtZj/hJDyIgtrmm9
RquLYJPDBlFF/rk9hR86GQISGmKk1LW4ku9PyIG9tArzZbLiKfvB2YeVqjAXYSo/gj12lgk7sMae
d15Yh2on6JfIPZq8JsWL5T5jpY7UBDYTelN2PQ83uU9pmOtRFZ/Ce4CsByYYamYxzo4xz0OvGH79
ixN/SRX6G83O6uvMo+PGvt3iUO4/j6yAPIBg8zYcqpjaBjbLueYzRyDKmuAwRYxaodCysYoN6k3j
YOvULU1bmlX6+V9a/1r5fGOGTctRJYQj5f49Ju1NSRhC6Xk+xw9UTooZUw9i8LkYc77c9s7soBOO
5rSjEnR+NfN+3hMtXEwFZIcCwscNAOjbIgDPYcucFs0pR1hMCt27WDdJbA0Lfl0PITnEUGURdVzB
ZKk9w3bWkbEGEL1G2b6ohGX+IpmBpg4Cg4hOeGdR3HTW8tCYjDhEQcTwhd84XKyAXAwak00CrUDk
2HZ9T8rIiQc8tnxJbBJUcCVYAIk+9FrebvQ5zDELQttM7QIEGc9ZdQ8GDwzjtQ2Jw6n/2zcbTioY
usK1rhiymtSQebAWblivQmgUmTR1Npvecz3DgCJbZoCELoAhV1SCVqGZF6qKAKiPN/zrJgWGEE7y
C11Z7u1FN/4rHvWCJ5LyDsxOJ1t8RSV+fpgx6BkHqJv9rm3RV0Qu3vHkompSZQ1iaRXzl//Y6FZS
K0R/N9EgxYYbpY0f4njEMXt+30k32DUFO708SuvSp+UXvDb3UtDSTH13s4iCYOTspNp6uU8ZMXrG
O9SsYBRWK/rJ/yuno2QnUzQ4aVzu6ZeVtaH1zEBE0xGjsf8qKfFmGUCMcFBx+oQ2ssa/UU1Wvqrr
QxZGAam+uwjmiVUe3/E8/AVtINpbl2zPG33wvdrlH+XW3w+2bYjkdfP2EhQX9rBfWB+mC046fYBw
pxrLsNwbDJkkEkRJBkXtjwiN/aHm5q7pAO7YaZbI65kOsFD2DGXLCnUt4G+02cxxG0ldow+d91R9
ghjaI2PoWWmF4Zn0tGKs63y9BCIB2b2Twm8085cFicxhTP477CMX1NieKjAx+Eabk9C76Nv2z6zL
nc04quuKJTeCgoh1vSHUH2ZHUTteVBsDuGXReTa3oJTwU298XDimXi71F//fSNfaFhn3GXHWIsEa
be4qoquUKxi4jjMKaX99x5Vwz0dQPSXgXC7JoZEmUbwGA0QW7PCvdlyE187hfNHXw8cAzTCIBgU4
Y7aonzsqB5EllXM5v6dG/StlFNfSyiu147MAobqRVWl1Vc9xKMgBl7Jwtf30O7rIpqQjM9cPLCwW
IP92SdvHBjkdMJ0Hkc0K7Aoi1JBKEAz61ld84k0MS/SnL6F4ouox6EaVQ6xY2dVjXdWysuRKoC38
xi6lOnVY4sAcb2ODJKvWMjYv5Rz3M89fWoaWxFcHGBblSgnv54H4lHAZ36x76jOkeuArlIpFqIxu
iAwuj7F2U5X9YxTODF6rldXCL8eZH56yMnexLiADu15l38WZ6E4qEfGRjS7rcOiZYadrrWHkb6iZ
DGV8fZJ1uEE+x0jyBAsmL2JmONBM9hHzfXfkduP3yplN2RgozTuw3XnEtkq1iVUwNLgfsEuoyzWO
gh8XDyVSmZ3T+QrqUZrxERym53MRBhaKrrdB4siYPYIbxM4gnvA2h4UKQBfCISjo2WXMFLEXK/ZP
+TS9961w2Z4Q1SNYlfuCnlgcjOz5hDvlesGVFT9qW5E09FtPWc/RvadvVwI+YEM9Y8kKbujxQsXV
3xlCPRbZD65pY87nFUlpYW2cd5G5azDquolbJSVBmaUDaPPQoqIGYYwXfBJDGY0mtdmwogxmUeSF
GTvawitHtZunS3+/XROhHgpSae8CMF9cAp+1NXuYLuNAVbiwJekY+SocM5/R7fC6g+2/BynXzpEN
VVywSl8nncYjttspZkbZ5pALogoyFxr8jGGxCHnCVOUNwlk5ykwv9E4uIGcePjPwR8/S5DV3CxkF
1GJGwpzP1qhKOXPRZpQCwSjefcjRg5Dy6CzTEWh7jvnfoqMcHPUCmAr6zADXiRVzahM1oa24MxSJ
KgSxOG+V+evWUbZ79VDIvM0PQFc2XqTTrKYJoQsOxoKZ9mlSeGqlMspATDl2E2WddV5P8Temx2pl
PhfTg3xAXZpTfWMJJJqeKMWm40bJ523CVgp7c4x+Oqm7Cs7j4IFwxW2Kc78AfAhUI30tYtvLBtHX
SXaQrc8+Hd0aqkD1xoidrokCbWWB97nD0y1MZJxFlpURMCxhTWAtT0qy+Np8iVh7SWkuLPa5bL3x
yeJCQt0P4XR24G5X9H9QVbtSqBEQ59CI8CqUvyypXo28EtXxPk7ZRgl/ZXwGcCxB1fQ9AJsvTQzS
gBcwUhCzDbJTPHKj1AS8t2NOz3IJE0qeS0Wx7/lMxUIG73fW2tgruJexexeDzxyxMCRpzhoHCs/V
9Tm6lknRBxt0yj9Bp0zh3nbF4SNEKNsSqM69hMhtBTLQ35vkh+OTLRLrTVMZPoyYCO0CHKS7lGbW
Er8BxFF1rLXCQoliXEVc16C1tfOhXZoEB4cfGQ8SMqMUFD9o0Z6YcQPX3XMNjdv5jFk58v5HpJS3
QHwphfuT27Y6x8J32pBOQfiklpDLKml0/wKb2OQ4uWr6vocce5P0A6ZWnMa979pv1/VfpakFsOWh
FeKFiBnJuBFuVOEaE7XYhU/tIDOPGa1JZ9/tjoSjkSvC8o9oQmjnNQ11SH2YQJGduP4/Z0bKAPN3
KQhqmxzYrW8ZIuyZwnQy1QTWfrcdyJ+j7RM1Gv1ygEM/9PWxbcsC9dAYDebs+1wvak9tvlm7kpyr
OZaKSpTD/IGCjXTBRoBUOoulX3eyRmVKy37Hd4dMUG/Wzn8DsmLwus0pJ+Q42Etz1K1PH267HQAs
bFlEF20K58vpjlTFu1LGT8d9Yre2/IQRZUVsKa++oP8I664MCcKoKJ/9BYDLNv1t5JDL10AIoJmo
XqvyVD3hRjW46WwoH2D/kbi49C9bE5JCGZ8l96ixprL1vyKEvETHKbuceIYlGOXmN/b0GUpFQ34B
465kjgOG6KPmMiekY4evTH5ELfpsySyP9tNwZQAjKFSdcoBd3zvLNjGVotmz7/jNszE/PaDhbZDg
PlKJdW4ZKZC/jD7exYZlgQGJ16Oz5Uub2PUXz9xvFk1rYYq2ZAJc9WUR8bIizxEymdQWDXwh/72J
qmzsvcf/uWJmQQNi2BcpiYdvzcRRF3RXK0sAU1V8XrYbA9BXrebDuHAae2Zpcd4QihfbQuF5Z6Pc
0yuoHdfe592jwYNzSFcZYExH+0wuaQgnnoKzbmlSYrrko3Y7MWOo3HytbgvksyaRX6dzuOeLf7hT
hvU8NS3p68SXWKJPQgmz/6rqFMTD3GCaduiNmAOXlInah7k2JPeUpBx1Adc+NJgjf4/pF1cwT040
shwjAHFA4J7WDkeYw8bblG5kZrEuiLPRRluGDeULgeBkUB04SUpxhXKBE24/uiLA6JInpVOZgbLL
bXHF6oDtYdSBRWbNL6fcdR4PVrxWNQTNTi254FYBkf1rG6+us2UQx92SA4p18CkiipbV2n/Jqat0
daCZ0drXtpFYqcnJkqQohe4+WTfOVP4PAln9YlVjiicmYpcGDgIrdAAojPgEfC6YLi2I+cJfzJHK
5fA4GZg7F+ouMSYCaEkRlcMCebO/+J/NfX/0RJJ5NwRshu+IQ2XzvuaMzHh3fDuzxgiREVOe0G6Z
ZLsEqIibh/lJwJoZmUKBwiuzLZk4ItGcK5m5qDKH1WXdlObEh6jQsW0P3k+mJwRnGNL9C01X10Gv
SCedLZYb34MXC2Q2h1qHqjAa0rlcDU+VUUJIVGqisNUCl5L2nL6yRbwt+7qOxg/r+D7L/iYbBkzH
xX5L0+i+4o+8LQOFEFUR0b9b91WxEWmEcPm2rIHwQrj1JCJER/vBTOlszRBJHL8JTRiSu9kTMxc9
pMFOIDT7eQIa1k/0EcinKaW9i5x/fR9mOaUPABr4zl3Fh9GNtmpZ/CV3x8QOo0juIoBEBSw5LiI5
XvWh/bmAsDfLTMe6mv4h8YgAE8PIJnVoSwSrDxz/5ttTqQiIqFeDuIkdbMilIKQbyz9KcslVIVZc
LSbIHyiy9Ww6quOycgGdSsaH7ZQvh9gOZgc/QzQu25Nb7zwg5qtmcBZbGKhInQeBDRHDVVZkR26c
7OAHBDS2wN9nT2qQN23w2bAGODtotdY1RpBLUds8IsuhtvHenM3QysAzF2M0LBUcu6EKoNGte49M
FxBUO/nAusDoDNgMPzUk2HSEP9hZueNja5o4hlkcOcEh1NXt9FtENDwbKZO5pIYdLllvxbg5vym4
lMZmC624pLJrXccIQu8uNPfUnKtGgiDqwijd9lXNzE5FDp9R53OtBUudRBOfo9PJOJoobg2pJFGQ
91Xl1RhCiF/Bw75fZ9IHZVwDmYx9zAbN7DflqGh++lDlDXQMxOf6GrFiPrXYfyOdXwS1OpD5iQGH
EO93zHPvLxBHwUKSXK7uAgdbf1qNLikTsdYjpiovZgXaKTXoQci36Ws3C+9gFeUcCJuqt9ph9OQN
1Q2Xn+ZWby81yEqJBz1Cg5jp6bV0KpnvXS16FNn7wEFDFoSsbjuZRr1AZ3WW4tc07KRANIzudgMm
dP/slxCht7J4GZvt4s/mIt3SFp4xrf6DSUO2V4CKD7YGx8nXuqqsKD6K141k12/144QkIBvJ9AOA
Oqtd149HAy+OW0kjSHKzVcjj8CwKNIhNujh/9szfFqz9rUuktXuE9ZsKm/i6V/cfJ0esYNrsLzUD
/NeriOqCiLkwYeeBZDfYnANE01wrXNKSp+e7TJYS1N59lhTxqsl0uQUpHl2gKWxXBQvBzwm3810a
s+I8bHr0oB2fFY9+e48k+Wlxseiy7avRdNT1aKu9yMrBrTqIWqmXE1VSwQT0ZONvflrXUbTU883U
kszNXj4V7sFQli7T+KAH4gSawgTYAoq39kjBNRsHcYRsfxKLUf41qR5NGpWiLZzu97dzdo+YJb47
K/Nsbe/g+ofF8q+jpXuPykPQRgh6Ds0wWAbfjI/srxk1mfygIrepF7pvMhnqg0FMnZH2SkwU4j8f
dP6g4tXtdV8yRhW+s0f52IMMpqmkDAEYh2fxSFxxHmkICwk13Iy+byOxhnvwwvFp+3bQNTRAGNyU
RANgxGD9a0HrIuEpYfgmzPq8YpgGcmQIOGIYKRVOWapBt5TcXaVypFw/aakgJDQ91jAfY3VhNuam
ABqWrodFxxJ8MsueQtr64qIPLZ1uiq0Cp3azVAT5qoOQP6yuZcJSVMVs8DajhFcvVKVp+YwJnk0T
9gWNTFwBbWwncTot/2NDRdYkpZ9rOX5C6x8yGY98J+AcRnHqMcf8wniFEw5R6+AVlPk2PRK2CD9z
ADnVCFfrhQs1KCg1pjO0fMkoWt64M3qnLgKhNC6Dk4yAlkCHjI0TLxX6XDtradZfv14DS4xTyH5+
aG3HXwLH5Jf5pCRQBBx72j8C3lStfqxL/rJolQIHdXi/yeePKv2UUNlnM/myrnowCMApKyIlzZPa
p/JMze3EZXg9wGJPzLNCVjl+xS+873/KDRj437AkNVXY60ubjrH/9mwJsrjFj+YHQWu/CkopkMBY
7Sqy8og5iEqheKI537NctLPFTwdGoRs+nNe3gib9736DeDRCo78lGAnmwjBYo9JpztPPK0Is2FLk
OnLe9II/t0K7EE8+0WMPzOF5rEboT5R6ZxQgptJ2wPNFURaacAfGv1IEuhiYm0vecb6XUAZnF+IE
tmHXpeYkBvoePGK8sbI/EtjsgKmJjJ9tsvVzbRdpXyv7IartFcuW8Q5OeE3OcgtQKVGEnqWJYAhj
bOCPLvk61qHS0G0LvpRi9X8+lQyF4+mGHYfNA4ls4jfr7iQV3vCgW5azYErgZQyaFLWrMNdRcaZK
aHWI5xRe1G2HiVnP283S3exBTYRaAC4/EwuL2t+s1GQCYS2ZSps5On5HHaj0WCzhC1d3O3wz01sP
+uElq72yJR45Q6wzFg7C/tSgmWyqspskAYc+RuQ2id83i7v9Yx3ChAiwKDL3NlTm4bEzQQyfH75F
HUvSoYO5vZocAdj9CoKxhjEmRkSV612/KKgc7f1aErpiUxM4OnhYUX8KJ9W/aaK4Im0fPqBj6X+L
gB82BySo4o9qD9a19/eH4fMwvEMmSrHqtttTK3QOKtHFMdj0Dmhpg0Q+lAWs0DyMLz2CPRSDFszn
Lb0f776PfgPlD//7hCZ/jm2SZjWok36kXC+oom0mwkV8w2L1Rh1jTAXj/Ds7Q6kfP0vKK0h1i4uj
JJAB5rKSNZ0zejfTZdXA4msIL4CVJIlT/ryB8KMy8alH01Nbe9DtV31z4dqP4W4fmVN/KrMxpiEE
aLFEV1shYK1Uw/O55ZthqxBMZvxsraWy0cLd7cn13zX7rga+JtJDl5cCLam8cdEBP3RmWmyqB2KG
qeop/dCVgpM2giDtQcnVcT/yHeCT/YKACtXR8FNy0QINUj0UA2VpV00IunmAjSG15UG5THHUFGC+
jeybbFMm1ptUnui82tFy4cCgvJgAzHu5zzknnqxJkYzHlEDyOdt6AmZ8ydZp/SQLZVngfqw6BdXN
7UnWqi11320w9ALS0j6TuFaFQtq31NDWcT040bbS5q3CM0WboBI81+kSmqs61TvdpT+y1OvSq98H
IzR/y12hndDJjFgypOFJCPq2F7No3BbT+yuE0Gz8M77kzN0eOWfcsYswHb7H4VBtXr9VvyJbtjLg
7yNbbHWPavWIBh1MBImSVKHG2NPI3YCMoQqbE9jKmJZxmSkYKiU7MPU1FGuz/fTY53BfWgIFUlHP
fuPsUvtkm1RgpU8r/esKmAueUFdos4sGHWzqtuL0LSgNnz6aoeSbZ15tFy1L0EkWijg3z56T2Rz8
ZZjvY/sBfXJQ4Pmy8YPWjSxSh0Mtp+mZAzQCvliUB+dNRlHZ0bh9iDgtyxYwDBKiRGDHA2SgNUJw
O9koiiNYYtk4toifWhQcp6dzhdqJ24j8nhGhu27oJKDxt1R/JwHsY/wSW21/SmsnHbx6RtVnXtUB
A3zByYgecVR3TfdnzWnqYtlVX1Ml1nylFB/IJCx8kM+/s0G4n4idr+J3bijnLc//rrjVHtnYh7t8
fpxPaC8ALlO64LlSk4/xd6WdBZfTJ/2y++Rg4JAT1lPEo9Ts7gmQAOJRD2u3qOVZUqzXG72ussCE
xXEDjtAzSTKmDyv2wrnDOzudTKKNCmh+c4YDjbiwk1j7V1QzfZ2r29/9Jwk9vQaCVZLo0SfPabHa
O9SPpTYrto6nJuvW7V6x52Hgmc6mTaQFw1CQ/Xdsj1+d7CIYJZAcEZyF3tteS5TcDzhlIJW8vcPf
9+JfDZY+kS2k4AQHUqFjYaGzxFJur48fxVQHxyogrQV29MYm7yu8IRJgM5D/LHsBaFuA18plWIqV
s506HA3y1PiFIyezAKhZaIUmtIrdVyb4nrQRVsBQlmYy10apEYSECoz3UnuYuBZ5ERxJzJnAUqO7
AQP5ytlvY6bbs6rRLMoQeJUpcnDacNpFUQWEhbTVU398i7h/AgXq+lUDRuxF0/zeM1aArep8BrKj
sVleNwsQhqYoo3sHWAntPBTu6Y9bwnQhGdpFBBkp1LUa+iFtqfQlVUjdrRSNKHwKLRMoYYzg+bZ0
KrZwV2sziqQMGDTOdGgkK0WusDlWTNL8F8KLnFiOqz6Xw1A6Mp7dl7IRfsD4ZLpn2wiJSRt3xmqj
ifLJgQPEX7DVIQkdoI/KAtm9IUCkdZ0dahHy+Uqbjy53LosV4r1f+n12fm3BIdEpHXxfHur4Q43g
P6Ohc2aBiinWkZALFfFARjQ7maVCCWmML9bxIdk6H5kFHRP5fB/dOuyfyF4cWbVTKbEYz63NWQkT
kxQ8OVPuZgxzWW6SYHB5ghHVRw1HFDUq6f5a3OV5Yy6Hdh+lKDuqQ4fQrZvOOFl5+xM153TaSiyf
PXC8tkKYK0ECPnJ9jHZgPRGXM/qPGuKmrhrn5Mr2Odr0LBLNBNpzaNwmAX6PMst1g8jgLhARvQk/
oph25c2c1mR6k9qKZy6HwaCRYrqZujD5bJHb2saIydfmDpeQ9G7ZHITOqN3ute2UhNZvB5ThKETa
sl9n7VbSn8wlztzn8IyV2JJocLiaJ4hc/PQuMq3uaRBoJeDWpDJ6suI8jux8BNA0LmmYqgDUMQvC
RVLt5zqtm+yWaYBrM+BWMhkhLdHn2VrB6f8UHAB2CjzqabKfMdrAcZevm/U4rJioaN8NV1s9uDiu
Z7ZhL7zXAjCpJZ7BSKY6Iu++m/NwFeUlhawrTXZRx4MeKAadH0u5qDrYCIS0c9YHwgeyWr30b59O
y+C2IicEWVdq7Em5OLf1NcXzBb4VMLlCihNAqNAxFzZAqnbtPE3PuvrxwE1NllG3B6ilxBOEZMzn
U9jjRLxIlD8HIyHFdauFwB86CiIzFWJTGn2eKiB7KNR7QkmVLi6QZz2NWKbmc+LCzQ4yVvgJSYcu
6AAcC8zuMJMgW9lr5oIrQSLrvuhzjg+YT/ueTsDhicVvXwyb2ywgClqfLn1nzcEbfioV1muWrqP+
zsBHXaEdS711YZwK3kLtyOTB/Ey1PASSyBwdGhmfg7A0WK5dO/ehSFPs/WeOMO4TdqLXB4fFxqt6
kANV7RWTqDNIDSkZuVCOOuQbvtqyoFcmAialPb4XsymN+ilwoCoG0kpYWMZV0jD4KiPDY21BLNWx
LafF2onQpc/95vfOmG+/4dKBwGb1GB6YdclLQ3VOh1yibpfzW8mW++OfLzKM/K9oH79Yw6LF+Z/6
fzJLTsaQVyP3OEHjDDLMAXYcHstmKN2QOwgMhplhfF0MhY996GyS+C4VjlX3/6YhH3XIzIhHHCu2
NzdwEITfmRum2AU+SW+ynfUoR2lDV7qnLRRXZOK4vKdoRmBTtoNYZ2S2OPAEPvVevisflf80pvcY
GqAXyKG5obQvsevYpFf7/ZTgioPynVcN0Gk2oAOH6AJAa530vwz7wn/pwtxATsrYwBQB+RhqwbJY
A3fmpqjfGM7/1wkXYzCkEh5m1OARFBPMIFLsu79+GzqeFBnA1F2ISwZiQV/UrHrkR9ca4fgzpbOP
mTXk2owDZQFBHOwrX201lcXlETrn0Oj5vPaUt2oNtU85pwYW+wje/GiKuBHHUzRH+DIkaqwrKH6X
Z6aoMWQdfn1BAgZpQYJGosxiZZuBDKAQhYdgGjUw/12YqUaTBGpm6VAAeFbSQoTfTtuOT98ZRDIo
LTcjjzxd0+ig8auxTdjMPyIOzEjCsT1xa9W2KAlErU2x+OV2QQNr4pv/atD3fnmOz+kzG6gr20Q+
7789H41Xi+Gy+3l+j5LrP1CnjpkhIeknjX+a+ki8cszUYoPoD2u505NB0E3/MCFp/4dvEkrd6cUa
SFZa703wi4K9KbceEa/qd3vE8RzkfKooWHOCEaXrJV8GjLO3Y39QZIU/PB4Tr00KoKYnQT8lprgP
UUXIpWfcjxXcYNVbDfqB4lWgINFX9BgNMpNdz9BAWDEtFo+9PpDFITT7g5IcM813fDH/RjiP4Chs
vhg65W+rYesldJnGufFaCD2zmWOMf51P96X001BmSN6UHR8VLwiPfccf1aK1IF9zD595M79uTRYj
l6TbgvbPwnp/R+OFSsAsz1B7VMwxBOdl8dJ5o8t0Q65xSpyFZjcppoh7R98LRIpQVKsCBQbB7Ira
sFr/YZkxG4p9CbCI/eLHAy83w5zVlKegjcfMFBg4/8JNIdi+zZ1YrTty3Mvk9PAyqqkDLlKkjQ0W
bdpLZROPqeYOra6PZ6MOqP/eLNaRbUlllrtud5tR44CH7AUFzIYnRlTt4kT5GMOmsmHAYnvW+7k6
ZlMp+bpQizB34vvdFnC6ngeNE/kfJc7x6kiY8EV3giM4lxfD8OhzrzLN1WaqZ5Jr4G5YA/UluGra
H2ov3vNEKEGPOZzLrZ99DMkroOQL9EcJNh7NrSK0yDZiYszyhr2g9fxOn1GTfhqI87pTKLc0K5aA
twWFy+jwe/p8xTzBvfPoHq6dzg1VdeY2CT2ltlrdOC8h5xU+PeR5BPqMA1FzaLLzZD6gD6RUZxOX
D9lgQMy6mC1ogitsznz4alHVG0oQVmqcm5TpFhcq+BAvT+b+vaLxW0rD7vgPgCu5fYn0BkjS/dlV
Ya0S6/u89mrWwWUbRbg6eWPtuSYHYYWHuWZFVhvIDKUTAunfJWWjAXqWQPJ9lCZQAG9dROQvMcJx
lo4fgQNXR1zPPqK3KJgnCNIWvniF5yHrminx+qFAFli7zBGuKHKrhfpoixSrHq3NuoNufOaOKOoB
ack8FYtRVrIItngGHzw+3LRnqr74w9q7sObV9mMGGEPEq8lLwsjFypgFC0QbST/M/yIVdPdmdcKb
oa+vq6uqv72crEie4p1nCxAiLI1TAdDg6Ab8IDo6IHOkc/IiIoqu7XiS9h3+zNbZzZkto349CirU
XVzEDvTAD9TpQpMnwOHUcz/mSjdRTrSlnalSCUPKM1wduAhkaBo/nxXMjYagPIhsGQ1MJBXbBO/O
RVYTOYPlodWfGP6JzNc0Iy3XMtAWL0hk9s/YTGN5EKdRuB0Bh9xHVlUv89hj6FWA5o7MPRFydfli
aBQG3zt9mHUBT5qISmBMWhEmS+njdUzHwiVzKNsjrNBqx+155LpcskyIRnnYSbi0zFy03SYmVjG2
z3bf/1ikwVr+Vu+c22wbHsUJYksjz2cFUQZl9XfLN60TXSbcjxidLX4HEB6Cm+1E70rTtNURx5+f
KKTNcejyJNHMyF2Eeu5ZfL3wnH9+OaO7g2cYsMJUfvi43M+UsiDGE64ZLptkQQcBpeD6x10XrGK0
BzKFE9+EzW0q2qps3DFBLaWNK7Vm3aVLvbnDlO0lmCGr2brYMi03vktDX9jnY0g8HQZTeBzBSbN4
gkOz8B5cvTLrxky8n0V/wLNdxJ7pEMymAgr1nANo7agiLpSoFyyY899lSIX1AqEv6syOJ95noNbJ
RVBoh7Ulgr4YSZbuzsCIb9DKts/h3ljxarNcmjKW6VLdxDEnIc5wt58DiOlj//XT/kwESd0naNXj
JZ6QYivjIeO7bD2zzeT0MFibGYYV+2wl8jDEnfUTAhAzQTTGRoxX12emBWZwR/PJKQ8vIQMVRUgz
B+TrJiHIblKfEOhZXFGE0EwRSXRmaPkwSqUhnRaXWVoRUkgcya0Ph6gzTFefUOSdHyrsx1bYKu7R
7GJuVRI5yl/De9w+jfAfUlm9r0M2L7OF9RgG86atuN2YFawURpGMZmFXFs+hMcMAQXFREyM/iDMi
FSOd32Cad09IRH6XKFHA/YgB6Cnzlu321o/TwDGdEu5DHGRIOydlGpwPaEh3RdwHAzFuFEFAZuj+
+YsTbm4Nj6hLQpICxZc5znSmMD5wNJC/WWPDcRnF+jnG/GvNey5WXfvBK/s21+K1WH0CYqc2mNah
6koOYDTaFZFDqVu+g2CkoCETKFD05XZj2YvOQ/bZthAacvxBxWY58DOnxn5OA/2LG/fCkxc3RqRl
LV6Z06h8KT/z/wBiNl5Zot7PBoU4crrfUw6csA6Tg7xjCtt+E6odFTwL5X3nzdpf9SokxvWam7OX
S+t27O/TvP+JeDTaJqKe5xo5RmER90gEIq2fLpsmYrjVP1R5bVcQ9WIriSUOPM05IWvAI4gK6Fv4
cEPpJQUwdTmT2ekgamebI44m6EsHaFqc4trrAuW38/8IyJ+64u+MmG/C35HTjnzIJ7bPda3OD0K/
jsOBz6S10AfTXKTH3p5Z5AOf6gl+czmnC3u10Ec1qCoPZq0sGEwEk7ayrk277+Ygj3Iv5XAOI7Jc
ijhJTp0aSDYUh3IFGO3Zu6cKAjvkvTV1tdaJxIJJ2HdRprMHjQds0sT8jf8PX6d4lisL2pcU9RgQ
O6ZkSp5P8OKTr7bWMs5OsozUQ2IeeBCYd3CQFjUkTwFw19KyCfBGNJFjd64kSs6ejYs+P6ByVOio
lRM3gQD42XdzUl6dEKlrgTfmk396V2hJdniduNPvdh3BzA3A2hiBWPVzzKjxDhpxTBnxR4jqCmdj
oaGZiR7avz+JDHbkvY1DwqhwQ16vaBxLAffA2++Pns64n4WDvv7eUlh/e/YsSS6ZKCzFEvPzFDtN
ZGRIc9L7vmH27OPDAi4giBhGA70SzvNx5MOy+7R1ImC82AOdkCzVqQeYMbsoHzvhMfpdnkRSBFHG
85wnEPKwQUi0prmNg/7q+KNmxEgqsy3n7n8AVX9sRthnlo51/5nqtFPJRDCfrCo0/oDFpYfVkZe4
hOG/W7qIpmJoyXnCbv0YU8aViWenLvzo9xandcCSV3fuwuOx6ZrYPtk6FjRiFZCNSZBFlHT2+YZi
ZDYBMhu/EVkl0k9L90ya14WRVivL383/OnIFJ70P54ODR1EiKtoJWs/l77Bk22xTkF6EajDuViBr
kBU7cs5PF0KCvV2+WfwCOADC2gx1vkjklPVR6KyX83rYqxDhHQ0MrasCVy8vviYDpQnRM2f1ZqhQ
YRpuOIq2dOxWQhKLuCimZIN5V0g7u1PhiEVSZwA2ZE/hJ+R10SRTopGK3t5SV6bxgXV9IC9cYE+a
3QboqhIBVXLNkjqvLLZ1u6JBprh+XVtBTnjVBjvht2VsuiyowyW0wxxAQAlGe3MmzJUN7bywVWRR
tRi2P9PfZsXEdK9uFVbjMSErROVcIZatEEYaLe5Z6ySnzVTBqAt+JJcbA+EQXIbPHPnZg4CXxzIR
2Yc6w+Lc/VTMjR0vmgFBvj4PH2eMfQvKZUXxYYYdeFqev9urbIEVRSIIMoAuRKv/2ya4tMIGk+6u
Bnx/Z8zDmh0rZYV79uRegs3wkl2VIE6lwzg2tLhaRX65FWwIC9jix7YlTbMWdOt1GWizpzLA9gSQ
Rj86SI/oaCkrByQ8LOyelnfOAFaJ8FbnPEKEzWxtFfxlDho+suEolJej+lKN9ofuSHSbnEJUvG9u
ZESR+3HNS7UiDJBFs6KF3xAqwUYaY1xknvopvV0iL40qttB+KJJX1Fdwj1NL/bn/Q3HMDZY7n+FZ
clQp90r0Gg2DCkJ0eycoQ2x2Kf87aRoiCxst0RF0AyaV3RihBO/GuQAKpimdkfa8Uoaxuab1FMcp
zW8AltNvPG9RWY0Q0x/go8HYJZqKOdKl7PyBZ7a9NXtDT1OS2Q7u6qcDh8QFYy37BWVqKPEi/8Ar
CO3M6oOrbRPedSN7+54qXi4aXAVoN0Qy3a1tQoQj4iToDoX21/6IkHMeIbklLSQl12lFgIPXrz+C
5nG+M+2x5mWE52NbouzlpCqM7s3pijIo3SlvFmPYtH9A7T79+NRI9ojxqJzF4EdqFm/csq5wlJv0
mBvONg2INF8bYVZlQW4X785z21QNYkYqR51JDIlxxzPZh0eGQFFyDjIofTi5oBSciKpDpbJ0C/OM
J//CKkViLP9TjGdk7dysTZbgil65D13QiBF++5Ld8dSo/nSRrC+vGxkWkXsG+MK3/ux4NdnXewfi
Uwg5Kl01uKdO++GAaAyr0rtHqOYqiY6V/jst3AiiF5maAwKMjnsgCcBQU74PFq+19jVPLd5xwMkh
iMe45Y2vCiWQGrDo2+VeOELPUVndWt2AVCB+wDC41ruJDWmgEX+tdRtsUAN6EKlnW8dOaVV0O5DP
xESV6CQb0GJKvhMrGAGP/k9MXlo81p7wEr/vSbQ0tj61AnlsHbWDRQnhhnqmmXjyA55yB2PwG9ZL
tI7NCqvWwOd57QL818XXCTzr0gQvpbgQatma98LqWAppsSPX8I+2Lr/Z94qFyEllFpkV26YBdKPl
x38gChLeLcprO2O+aow5IV/eCCKg+9pN1//1kgR2Gs8L+5hvkcnwF3MYCNjYlnvyPf9BftJf+WYJ
FZuKMqwcjHTjvJMwp6L2gCHtbYKwvf07uVwZC3Co7o3vThF2UiEcM85l3EHK+7rbuz+aNvvDOn7h
7IUBc0Y3RIGHl0SDXJ7lP57pMgv9IOPRQx9avv3Hssc/4N9oo1cnv7oPXJ9lJnvXZWDoMgDjeCuN
M+9PIHsZijySC780wWgJ8kou0x5DVz3Zm0nuXIBaMfJ0esuuvqb9RDlmSYxD9ePa6is9Duz8Lcw0
ZtT+6zeb6Rn5S6vSOGltBpDaOemIzvVUme/Rka2soQpP4q71MO8/nVqdx6rZ3P+fIb0rYep1Rfzz
R2QTkZwiCa7vtaAFErYTvcwlxRSpgS9elZu3XC0OuuzMKzrOY7iHJ8HjtSNUvvYHfjVRsAfjOUGi
RY/j26OxixKJNXnwK7rEFzYewHO/FXTxkCe6g37+W1WrMve+XAhqT5M92cqVzmzotyzFkp+ZzV/z
iUjNhIDLIEMdrQZ/XjEBlYw/rj5xXWwcbcaQwb+jJqRrUEyFH5UKQJY5BsGU41lFi3RXZX/sM3BO
TWIMJe4rCf6Tscfv4PZiywug7wnYcXGxEvIDf1u9WLCDwAa/ht5JPKP2eo9YPBYcrquUdz9+iGr8
guW0Em6HieMSZRLfvBhzvtLK++93vW7kkVhdpzE0wEKR976tWMJ3xhefzURiVDO6EHhqN3sNMPkn
figTRwCvmcKNkQf+BTzRRv+Lq2vA23OQDGdxvXo9r1CZXhgh4gKZYwQRnuNXqZ/iJjbR1VH5FEnS
w4XNnzTop72Pxv/NCsS9RE82JgeSrp+uMQ5Mk72MvwbiAl/q4GOU3kQ3vh4dOqnkKwjbitJOxBPt
LUgJPIFlXQqJV8HNP/xphXhmKJUjz617b5Fv/NZdeAQPexp1OTspl1DwLpqgKO/YMhZayhZmw6gI
y0nNEW6oTrvxQGjA1Kv/gT+tqfNCQHNODcxbkXNStns3dUqHhXEyaR0SQqwM175x2vdh+WG/od3q
ZSeoyicIoMXv6Mx+1hQXST1A4rg0HHinylE5CdeQODrOduOult3NADKFaYNrKzfx+RzFfznnyG84
Yx1XoEnsyFS2r+M/qG/7SjKd6XMfkdlh83Kr+ivVR8/A/ADbtpSLYyDRLLTFyEZCkMH7IwC20lss
8R4ZqDc4KfFt6Klt4SV4Jh0LgznhZWMuvY8Zg53Dp//ujQg2jc13+11XbUD58PtQWu6rDbzHSVCy
PZM35RYs13w9dwdsjlSQ0yU2dZlowyAZpPy9RlldX/QB8HtZTVRxPJhmmCL11CmCJ+dQ3Zz/tITe
D0Rb56nD3V07Tw7Nad6iNCvXAWJLg+Xv8rVUfJE9PyXF6ygq7EOJ1GaZ7WwbPIXwnWjDb8IR87kX
rZYvctHT53Hybr3MqkpFU0i3sQZAO9jFfQdZ7Kok+lw3emDJ/xDQdXIXa3bcQbKFZQtdYQE3k225
DQEuNpMG1UgHpzk1O2kobF73aK+mLFOQ3PkowCxecNlJyFom2OMcUbWIf8ctQIK2VBCXU2MDulNx
93erhxmSYmF5PIjk21mBQTHvdNam4wcw9kzd3IHUHSF7qm5ZaHtekehIxiR4DcOq/xRYx9NIiMd8
Nftbw015vyFQbm16MMWXDMk8q5rkP9RMI7bnd8FWl3wSrjiV7Y6/bnkVjTHxz56IaIlr8va9D7eH
PPZ2w3SODXKtOXj95gJoAIxDe4phACKWzAxoBWX/JlOwD9j3ZDS7lcgV+6Fzsyl5bowva3pw+s5K
h7CHjYdeXCADFMQQMuDnrIkOCEQ3sJcbBe8JBDsKQuyUglLq4lG54/NGRycUF2McU7qAJKCbMIX5
dBQyl2R399mLl9qXqgd6bavD+jb2oGlRtXhvH68x2UcdiFKXV1LMuu7BbAGPMClPPIs8wMAX4cfV
MJtJ+4hGG5KmuvD2Mm6r+6kuYbTFIThL0M3Rub0rrM95JKOuIx/gcHrHdiHQQHSrof2vVtQz9v3V
BKO13aIZxmqhP2qSEAKxZZK9HI0rPn9AOr8ud7xCheE9F5gx7rkmKW0MZMJVE5g+ucvR2NDXcOjl
3W8qIy9NslJeRt3tjhDBA1kkZAZBt1yoRhwO2appzVtBYEacJSr8SwEB7efOPgY5m+4VbWTKqb2k
5Nz/0fvetiwkCUD/g9f5zOljw5QMEsUmrDtM+d+QLFrS1VZIcCBLkZ/hkY2hxwn9/SiffY0nFUl2
px2U0WbrAgzeYfSd35ACfffQOzsux5Wj1JO5CBW+qvPUelXK5oDUD3H8k2d2Yp+2Atymct2kJiDv
Rr4Z0b7MOjlCj96WOfeTcj+S78EBK2PsqwQoSuUO4GY0HsB4PRoTX/TjXWFiR8s6Bw/1CsWkWbc/
wiiFvRN0NrjAnllkWu5az/hZxeNG450EKStBzv9UQg1u/mL5VeMo4wNLVez6fytjERgWxVbN0Byb
m1I2D/b1WQ1+xFQVbR+pErfcOJEGwzFa46g49H8KgaB/rPl8qOSK81ASuNyx5uvx+PJHPntMQMsL
COqj5q3MYY1MaF0FHf2/SUXxJbKFwxXlVrzFti9G/Nny5F/i+iZSnd7+w4tsY8/m/tpf/J/Yru03
I3nFjisnUdjzcFg0St7Zjjmyj9KkZ/Tw04p6QBVhcolql78EQpih2Iad1446ckFqYMatO+RxMGNT
N2/gBWncLDXIZTSLu3bWboPglQmZoxzJk1ExIp7UfCOWhaWN+1VygDAIGMw1XorN3yUkb5Mnngt8
UyfurLtWUz6UOdP2Fk6TdT2/yIYjcP5Qc9evqwbLyik3Ce2CX5URhdxvhrXu4VYRQiwGsWTw5of3
8rucAMqUmblidVQDn2tYiBKxE+5GYBWZeRtcBDSaQ8ZXEghLCQKB2uE/4t+dNEjYLWoanxMqjmlD
fKNIzI4kY3pkBrHnbQOWQBYW/0Oyp1dfFptQlZM4LYVYG0Nluh1/cFMiMqAwIv42PQEpImKiUXL4
WPWIOo3p69z5gcUphWH9/qVhQ5GIWOD00scSfsgXURcBhy59NFyFNeSrYDM8PmrmungnTzVeYeLx
8GfEqNd0VLWFDxpMpffabQP5zwiuUSmGM9HQqazwwjZkuNo92y7r7vxn+7rWn6HHYY741XyC6zfI
gh3CJPVu+OO5IxhvFYtap/5Ucq0eZalfWPBATVXMugRFKQ1mSDQvm1Rltrz7UPgBXJPiM5Owjaux
ebJNvw0c+JF9+FDzzMVCtnetq8YuEP991b0UGxX9Iw4Vegbc1xBWS72fRXdXe5DgRBDOJaaidPLc
SvgF+VJ2ATG5bwH826BfGYH+JVaiwRtPBwx471C5XHr6Z6U5qRSsinG24w39wzB29v77TFoSDCEF
TT+XLboTfdFH90xmNs7hFz4HxSOYZnFgqqVNeuTDDUo7UBlzummXG/2IsQtTqkG4Nh01N9yo1gXR
m2jKCgpNfWif5JHSDd+van2Z/acG4UBvr94MeMFYn+49VedSLKs517SzNqSD00tBJj63vsTieRnS
XLWKPU73NTiKlhKx0bpTSOxXjjeTTBKOxnVQKsOaRLB6CWIdz0S7bBE7xYipSGjzJCjyXRU+Gq/H
hmVmPHbehJLmNe6c/yqANb6FlozQ01+QRMNIjudVL3HKL1IGFrL4YKvUR4FcPxr7kmsliuYCdYSm
rsvsGH9vD0PVH7AZd5zxX0NMeNkk/HhZ6P7uH3p9eKjeEXWae1b4k2VPifL4dvlPDdeMt+2Oi+PD
IkisRURFRDLbLX1XsOWz9R8xgJvK34+o0pows0+ynRIZdCzjLegptfg8r2knId+eBlGTkDx4+JFm
m1Hh23+uRKRw0gGnEcRXXJicHivxWeMoiRZEtq3YcQhdcSREy9BHOMvaEF5xIS5lNsVBKANeVIjz
VYk2mZQPJE7dNXKxPUYN+P9tGZ7/jpAligyxhOKP1gvaZ8Nx3ip/0SnxPyEpiiLFS80yxEq3fkIL
ymxLbNtTkG7lpSKfUO1xwwy5iSZ1fxqxsQOjNvX/uYu6LXHq3DdrIbb6yAdRRVPtDTr8D3LlB78Y
xCJY/ARgBAWZz5DJRdg4+hwJ7q0toozUJzD4Rkm8iNzjI3HsmbzlLWgbMlo/2PSsugaqkroI5j2S
OQiIdll2O5elh3uVdmjJUNwTq7rekEROPhwyUjrXhnqoy+/qnktHH+a736pcmFRVImKXgwec45Wt
BXijwScN89elJiwfVgB78OFKn/NGST09rmrOgBsCA2JJTb7LXRxbh9th17zsj4BK3KloPSIeajQ2
PHLu+xFYz+sWt7gFKyLbM0dy8oYCWDude5easO1cfkQXBNuKiw+GWOl6qNRqz7MN5Nbso/aSQKNF
wq0uy1rdwKaMh7COc1ayPQkfyVUwPogPOhuGvK2f7JKBo48FZ9s3VWKxhQL35ji1pyhJwmYWNsOP
9hIEodkOVTyo3e4beJbNzRSuqmV7gBOOfcB60o0isU6iGWYsUuyAkIi/Rzki0RJZKNN376+5lTu+
VmoDF7wi7UlcSQBS5tut1TXMP/H77mbw1Ip9NAWYRb3tKcCwbcMxfQ9iRP1ai+Xl6IEkDmYJE8xg
auRiABw2Zoj6sUEQmvirF9NPV3wPvVaiiA0h6lKLf+ndL814AZGwoFjYcUuIXA/njsBzmzGXPQBr
rs3BWDqXZWRRU6hW92Uk56s/lQL1KnGGPGuy+6/Z1Xx1lzji+CX91Ykrp8Ux6InipN0J9X+x/nKx
JjqbYueZtUEb/Vo/LyZvt0kiKQ7XEFxK9UDidlgwdq9nOpy8XJcv+fxIBgIA2SX1GAR2Cx0SJ6Sl
8yuhICmRhkwDYPWUUpn9MkOfqPmvpVwy11ZBVjHMRR1SfyOm0M546LyFWuL26v8sT15u32q0n4ey
RnrF3chsegoOcRUsQc70TR6ySw1PeaBWADYiYWdKxpXif3/m6meDZm98lulzX/dBAJruS1xGcHRJ
Xsnh7GkSovSR/LT5QDoZ3k3o7V7sY5+HPt/TE1G7HFzlHqwJSmhmRcVB9HYOEOXJ4s1DezV01ngV
QAielWfkobNkmL2YFzHmM2gd2tNE+K7gXPgcBwG9Zv/RgNm9v0vesJf5GrgrF9wERcH3tbSJtmho
rMfiJQlhsDqHZuBW7rJ37h23Bahb0dUS4Z2R9s+b98oDWWHy1+hUddAR68vAf4ct9A9v32g0MSDf
nrw29QVNGl+geBQVgs74ek9tCfY6IeDJIFmaS9KfsKlF/FU0EZR7wCYjfp4vjDvcPT0JwiOg3zIi
rIQlqDZnJLDGzvNuhx6BFZbyoLJiqOlv7je5lwQu9Ec01UM2q4izqQK6/uLgo1I73jAXhPMm0GHs
exYVB+6KpQkQ+/+AuQCU7gmXz1A3MEtpei85UFUyIMnamue/GF3oJE1kKW6i4oUcz3l/riYBd8uH
0FZ4CSjtSkXQeCuXi9XrR8WETrBKuuU/WvV8MD6xykH0MiAbjv47ME0VSn4hZS3PJirZ8qBRYe/a
1p3Vn5po4mLSlczlOcc75h2NIc+oeb5RTqaakEqzyE4tlEzVLpmEVA9tbGfH1RjorzHcBRgDo2e3
/o42TIQ38n/l/S2RLg3jVUeDU/e5G/jY98PwmnceHgc3bQrh8n1AYxr8ds1UROB1Yrfwx5IZ0VB5
qpKgNtMAeCRcVyW+HDMzSxO35ylPLt5+1vrG8ax02sY5QVc9lB2PWhTPn/1ruqa8efJ5bgmAcFLU
YMOW0qS3Gm9IzQUz/5++APwWugS0plwkpBETRz57FKNc3BOGeaDHcCMsAH37KX8RROu+IuzKNiWr
JCbISNI0JfyPOFqwsBZ/N5UrItcviLr20jOACOe7wsTzuF9jAp81mklSqBARZIF0Xq35hluXbrQC
jXM6PNlAhst/DZ5le7ZHtCoCDWN3BntcxspqF136s3LNufbxQjpe03HWZ2NsCXy6PmaOqUnFNTBG
kABOEbKrgKohmby1VYmDmN62U36Q4egl6EVZotE0SbgGuOfO2325tX2z16J7wCc7UG264Qi3F4yU
WD4ZKktnttc1i5FPLRjMVdqgKkY6qr6LTJux9BKcZQWhjpyFC0muZ4CsOtkXYhGF/aye9PN1ruFp
POO6wv5Cjs8pK/q/Q0Cy0Bbh4SqJL+eKVG+39DD2949iuPeY+sSYZAHP231mrXIyxUJLGyxNIXhL
Uo+CcZxq/lHwd8St4GkEVV3FEfy4tf11NPyFwi/OuDlwO7MzruWpWmlB8WI/DjHZ66X2CwdKHx33
vLs2BgrbQQCHSa/4I0Air/yCOTkMuYvtYv7YKgDY2d2xxtoNV/lgDvWA2OuMxxLKZWlH4WTQI6q7
3859DjU2tDIKnAU5NgPgPEY8yJcQIGX6ZrE1LTZCcx/x5g4alX2DnI85vElNMxWMfxz1NfiqL4id
PS7PVJFjMpFJKiHrtb5qLlBIZx8m7ZPjW1sEZaCRHwzKSFz9ybeln9kOs4e87IA4RBRWaQPPg82T
KmTb86LXwOZOH2bdhcKyhoCzS8KEMyqf2iu45BGVrCdbdY9yZ18x5eVph/VJWt6Jm1Fe0c8J6Vim
Qk/XLJHdagY5K6eXWGQNudG/xOIBnd3ah1EiGnTqcJHJHbCULjkNK0YblkiIWMCdA7BHeegzRZ+L
ASIt3FBtvfRlY/Lu28hhFWOJgT5vZNWvc5l99kF5N8+xJ+dpUFRBzHU3S3TtBr4GJV6fXEtXPufm
xsLhV7fHmqZJiRmK9OQOC7tSAs1V5r9sPuvLPI8bWOMeS5ikpi3TEs+1hDkSYwW0tIAIP5XXhnxo
yNpMCluc7CwdDqyj9MYgV86ZddK2eZueDHFNqUjy6nVmNG23CuA7jW9EG17VR1eKU/E+THBYQp8o
LCRKgcHA7sIYrgQq5TSCsKC2aecV6Pyw9WWaitqw/hmT8iT54VFJKtdtu9WUqLHmA7rtt5G+ewLE
zkAc2pOJKLWTiNrV2r9XmiXv2G+Q6tMMz/RHn50PkybX034oXjux12H/8BMOclMPMFbTU5ZZz43H
xi2w7nhOSQ9yVy76Z8FHFU7xLyXdZe1ohQJLGV9XNqueBdHsEtOQZRwBA9MgCiri4LsfMRWdxrSG
3O8NkJ51jMOFcm4mECgHe4TgIiMsvj8yzsezz9jSuHgt2POcTwvpKta+OYPS2G8Hq3QKgUExCMOA
EPjiFKo/RorZo6EkdSFeNsUG/92nrCF7uqT0moctH0hT5h97zR6rgI/HrA2OodX+YR+Lm74oLPJd
BtqoVQQNNUHM6BA2JNuauqJaBCspZTiWdL6IGq/RLgydNrMnhznqT8wgtMM9+UTJeG/ClWOiaW6J
lrkQDEUciCtUdNOyYnhLVRMTbSg/kYwGi2l1m2seFQwH92HS+8Cmv2OTnptB8grAVp73hsQ5m4ZN
qyPy8+ddlQxwTZMSFknc+sN8heauSiks9iUzDK3FLI2mJlgRmhIaNIOFw86z56NMhQ3nyMr2R9PC
Kex1rRA7MgUJTB2HuQahWxtlv3SgwhxhxKfp4dqJV2EXgQZIZCRTEdUU/e5neplnES6YepeIfUzf
7I4ex5kj2GXINI8jhRRgjT/jhyWuDYn21ULkk68Q9XdrcMn3jvgvwUt88+q5next3UVI4SCSZNWz
BvRL/LjUVPpYhnty/U50r+DcZ58yOBhrZLUzrn+E2yxygXpX42/o5pZekbMXAahWHD7zsf/Fu9c0
k8Xgqd72xPd+DVrt6GEOByLFQjck8fGAxsSrSni1uCKuhy/xuqeMDdjn0oi+v8rbUzSqGHFtC7lD
y73UCo8dXbn3SKKlwY1LU7UfCBu+LmtHxK/Gcp4w7rn2Io46+qNRrcAQ6ve43iIuwjKxlJdPFe/5
cj9xMdRkGld5MF6A2Z+imQlCgib7+9Vj1VZN9mPDqIinOny7yqjERlMk8sq8P27N2iE8KKA/nJUU
Qjs1+9c0xIL8EMJqZhuEpYRy/nxrOWH3dGEk7EAPpDSr0AaiUSjr8MtGzPuUODUzyhyGChI6umSV
dkcM+pgj3Rs6cxtU4s2xY45tfeVjc4P4l63BVbvuvqeQbkoLHHLelbW59jrBGqutvazZy11uZzNf
gX9rn9Ygaz3bcO4j9bggv6ho2HgVQh6rpFwenMAB2JR26yzblU1cHyVRyVQOe6EZYIBzHMN5+KZz
TD1CMEsYS1D+v3ASnCcP+OvtS4K6GK1MaqETdA/mH0CfUQeG2KoY15DedqFdW8KXvEvNif45Lf0w
jUuh5UpR0Dla+EdNQym1ghp4BZJMata9d+sCIZh3/o4rMxYyYedCE+p05sEKfECzVed01SB8tQJN
9YoEaMfi+HZtRD+4D0ObD38zHqalRs/KlVTd97dCSpJGvvJIUsjP+aiWL+7KkLEk6qip83hiD5Wx
hLNVkyN6zT8m8nxHLqCNpkOHMMmtClbQCnf+nQ8a2ylio+7/cR6LYFS1FGvEgjjXlPMmGwC0u7Wv
y4zLU+IxTSjFh9zssNc+6vQKARed2HA/I+WopEvRnEw1H6+8oNFdbkElg83T6JiRbO0pJVV60RgY
QrNWNmupfZlXn47xJsSHa0s2bzi41fVG+1tSSkuykDPsSTdN2GyCHq1i18uRB+63YtT7xjlUJ6U7
NZ+ELU7Ph/dkMP9DCW5uEHa/Fe0IXxuOyldA+pysimmtQScATUjTe7RmWQe/a42gkqbTRsSSyyMM
SUhNdz6wL4ZXb5Lo7XFsOlEpTTXkns5/8hpVQj68UjKbW3zkQHPMy3eOCKUJ9qIhtrQwJAsw048T
0kFUjvuo/DC6jxs/aJrdWqCBNpQtPvzCUvtTPpJebuVbzDWLCBWO7c8b1QyQ5njuBOfxrFc2VPXr
7hjcdQz/mbnBcXUfutIGUoIDybnB0d3hsvcEBmdpS7WNUA/FHI0CBfW1YElFEiplq+7lRMAaiL9c
MyAKbccsa2ChhI9xm2O9H1WJaLRol2VPMqkIahCnoi9u02Io0AUwji42UmeKe6+L3tsnI7+Q+SGX
BYJZbQE/8nf7jZCosvbylZ38kBb99Byxl4Ii7680xaekc8IWNVkdQ61JxkH1na6UUU6y43EHTHDE
i/Hxj5iT5Vcz11QNbtfJrn76GaAL02j3kSdOS2P6v6j2+ecMTLS1HIjSramuerR0dbRnqg20bo2/
B8+kO15AHemXUp66D6hIn+Uo/XwUTtW4QCAXfP+vLCJA07u90NeABpkXVz5467O8gUFj3XlZ+cR4
YAv0Y9lxTfq+HPNZjuDt9PWIFnGPIuxiiGeowNpHzYIdT9ctYBkcrgdfZn8fU4pgZbJWgr5lgLra
InjxeXUl6Y2usMHRzeYDxyVoe/IkZ3dy1IUeyHOky8zr/JFFhej5e0y4TEdwC8bCyv/olBaZSq9m
qdI+1brRiQs4wbVKN9R+DOEJDXfrFzHyljQA77Sh5UcoLYijonDBCgX2Q4juIfNzOLjrqJLL6yzZ
iIwy73+SWl9ACMO5zo/Wun5B+7q/AD4wvOjg+F38Mcxj0nRctNjfN/Vojf41woLnY8XBcrijcidL
aCnh8I/oKFLDyC9grwi3SFb1KegA0tU8uDer1HTeKj2/lwEJZ/4TN1GGEYT7kG8aCCu8UihFOWOk
VyUB+2a8ooSyC19w0q2AKAh5J2is1zfYtVI8ZAk1145tGYCePX3THf3Wj8rcNwTZCyGlEz21+LSt
J+MusQuaZVRCIYYNk6P/kz5aiafcNYKjHAwEX96Yq76ONDIT8sJe7QNjoe8JqNtP9rcbVczT9uI0
PeCBM/OAMdvbQyTRMyrtqabqrqo2KZKzodC5BzLlfJ9NqLf2e3TDLaP2sevp71myMLCGxxumoesY
O+XP8qW32ICPQ1kEO9FKLPxa6ZynN/UB+NM6czqNjsOF96jqkREql0TgaWTUyVuEr8CRF5NhOXv9
EafvAwA5csmknQjjgIuGKzbotXq9sm4eIUGw7Uyi2XpYdY1PpncuKCqE+XqpSwfJUFy1wkBfpnkm
1RiwzfV6EFwMk7FYsX1+cLqPT5/8UvGVCeiZ2TBhWVVr9FaXdRaqKNePabynN92SnJImKRj+SbYu
JipMlOccPgtJKBg1M4/ZTkNBmhd1YA9ddHYKGi8rTKNBhT0/d7kv2vAVn9VwCVzeuYmlpPESWmVQ
67nYEuI1lkrJrvazZNleulNLe335HUF+5kqoe4N3FyiRDwri4by7H6anJgFgEUSpHFzQNVMYw9xL
udyJ0qm2txh2eDJcL6q+iOp+fZer1j1SH09ZVkDmoAhyQgxZpOU89+qlPxY30cFMIBkefRFOSMJA
x9mVyDPfOG48cXMDkwPLgbbSR5NWIXjuz75w17LL2CBD0Vk7LexYPt1M/McngUZLKth5sXxlc887
5DcVv34bNxq1z1ki5HiPCvdQinePrVLNyq2cRsUMcsG8TZWIgOTAw3pY6QA7K24ctW+TLDoC+VoH
BQNE61zdwQbX/vodtABGwFkWWPTkSfrn2T25r/19mO7v16h9Do40dFcFAvZbOMvSc7Tas+xYbBnt
nvOG5CrFeo6DEavVt++lA4aOFpfkU3WCGaGAXcAiQ6PKhc9zTdQLaG9pAOwwQpEZUyEgVgf8EdJL
SprMtSft2Uqa0Igga1KWQN0H6dkxxnHAVZPLw4PJpk9MXUmNG2gU1AMO8GUZwI/T8XeYXHQraD2e
fS30EFZD14Wd+/lJ0w5KpX6aODg4Bp9P4/rcSLx0AOkC59FqGN9cSqYVb9vgCClgr0yCR84y0x7J
6xNvFsaR8IUe97xybbc1b+8U0qc2MKytnkTlsh/TP7g7WC+KDFlQTO5XWLwbUNMIUMonLTcMFPFc
fsz2fJP1RpB+mOgD3w9+4KPn8CFwJNGae3ZyfTD48UBI0jWD5eNiu3hwvRJeCuo9fa54oTqBQQJ3
KzOPsHynwVCp6mbC/5e/Iyu1tQEsJWXtr0F7Q289iN4nnRI5SD15kCI/SsgBPwxzzLO+ByLS5AAw
W/oc4DDs3we1bYPtdgKo9QiO3+gvxr/AkVZTPlE2+5tNy0DbD4oSsp2YVSv4B2NubNfmRtquRbXt
OK6zUw3ssdd/Cg8NkVKUbj1rbDpWpHY7MV1txOJhnjSdO04WJQkm1sCN/WwDuA9cJ8jiBIYi5wsT
j1Dr6aj6nCpW8Njiy+8CLBxfXzuinUsKEY3xJFb6OWWylTAYfIclfM8IhCQLcltjrSEDXjf4Nsth
R6tPgscIdnOSWcTAO8EgRUrVdQ+JIRawznpJGJsaVL+Itlx+x5XI21smNTGzBuPj3QtQkQtFCNRm
vDrucnzRHkAlQ1ri6/h91TTB4GNNTfHLplPeIwW/h+mEik1BSmOYAJPLjjJ8QHdVR5jS4HV+06UI
+zC2V61hIEsD2NcpkXsVTfZ41OJjKCeICNa2/ImyGTB4EMfdDCSeWjIP2X1H9YHBd2+VbndpOgeU
kxHYD7HVYdobdaFDcLV2E9HykKzbAr2k+bnJM48/5JdroZ9BNccoaacGITzuxVoBbm/ZCaAaAlvh
I0BiwpRCGu4BeIHSm1qWux8TIavI6iJ3ToQiYnhBjYqjHZWnZ5gL+TCNEopY7VGVlLTQXfirqW8D
LmZwLWtxDdCu5BQF5O7qIzoFPEonxSA5wUHFgEefDIex7AL8uo9hg4GpEKYXXL+5S1zIwl5bOAp9
SH+qnfkqTmjIxraZ4h6kHl+ybTFkho6ZMDS16ZD7BhUhLEWCVwzCF/O5V8bRG/g80XWyGds/FXZg
ixmR3yJ65fVOisbX0IhSkst/fAMRBGS/5S7HpdZ+rXWAMI6F1wAr0LNcQe60TBJVz2Oz2pVOb05D
/R60ETPq7LHoasBX6emg9AkEPNeIbRm0cpC+PWsuxZi5jLmfNGxuPP0nMWoFwcdRW0aGWE2wKzn3
UgCbZ41TrUIr5YBMden3cTpeb7f64AlA9LZJ0LyU0COys762w1RCfTbZZwI8mknEP97K8AfVurBo
vwWswrWnh5ZPMxIGF+0Of4Cg7hUSajfkk+BgTd2eG23uOOkuwG0SErXpVGkG/HOygV8jFbrOOzxQ
p8MlBtBEOpjUZtg8YSbpye2p8xY1wRw62JKha+xPptgqUyQCzU7xT6TaUoizuBw8jCt3ogsAaLPH
tyMTODId7qgII7WK0iSAU1DLV0gE9hyOh2L+tIfXSDqXvSBdQm9rzdAPs0+Yxuz+D5xcmyfCooCy
8CyjxLFY/IYiIGHG0ShnA+Xdk9Fa6kxk9b2yPjb3AbB3OR/vFUFpPFWJpPvpYH1UVQx4/T8rwgVr
nrp1YvUJVyqbd686LIwjeY3rvjIwAWsQknTL5LK7D7cCb49FkMB6Hw1syhOlE/o40Q+lE6Mzkhoc
SAOUS9coPyjTuQ59pqYBM7N1ufzC5JdwRVuo14gvKJUJubC3aAbtGrYQI/hs5fTcx2Mfovmu4Tn3
Rdfakw2rq5DmGjw62dJYAQu4QHL8JpHY030h1e+cQI75/8n4cH9uIG48C+cmkaFm+waIAzekwxKN
VFdLtZ/yUQtJrOgj+XuVkBGcuZYr+iodJAKRkAaGAmx9wq7BQmzanzi9WoR0CtdyYjibef3DLPu4
kjgdBmT67T5njmJFmAUk/y9QIdbPWtmndTDwakP09n4tIuus/RKN2zA1t4rVqfrx1o7AwWrmGcy+
HVhKdiqaxkCg0JKp7HihTP4R84YNMW/zMmPgMGMTyZxYl8+MVjJhHOVinQrOU4LwEDN0vZsf71c3
ukGxgQ5FIhh9ljVlrOepoFstSJuDxuuGNAEZaWnbzV6GElgyxjbcPRCmzY5zDMZ9SuBkWWCzdPHn
6NhlpqFIkfl6fFqJTnmVRAXQfusC0A5SHLRywWJ1ujPULmjyPmg3v199E4/5GpckVhtgA2HlMYI7
x245hveH08kJ0AwBV+0WFMyz+PAAtPcl4ulgL8NAXLync7wU+HZJgXmhMEliCGZTC73dQavmG9aN
KJ8QfCTqxM1xxddLggCY/TejBcRhxt6W+zwvD7Y/YDCMf24gdpW9/qwv7usF8YzSMiQ4B+vtJb49
CA7+DH4B2jmdPutd93YXUseAzR/099qn8Grctk4QUEIL4MifJgAEz7rL5QpxnteBjFLCvuDUvzTS
me0WVd+gBHzcG+vH4VAfagFwBJ/fbbgDSGZc96fg/A+lSHP1Ibmw+xNfdSp0s2sDVrQfIWbLnUFm
7dVFTFNKqRxta5NWLbt/Q5jUDJTLWQRSlcZjoVyA6lBo35oLFEf5QCcEpEGbTSTw/ngPUeBEnBv/
xNO9aNlJgpGBAfFvP80eMu42S38pOeeiq9PVVR4uv97p1Re7FfcFsvvMsns2D9iFJRrYlfoW9raT
zv3ydAkIIap8LFx7vnVxlET2AhyGCB8UQzD0zg6DMVPAKUVabuNReB4NiCSh0IVBBwEsIlK5KpH2
LxN+k0zbco/vAHBxl7ok/09+Fqm0BTGMdQDGRYQN/6VbsguZseyjTnF96r0ZP9VNyp1xHgYzqanZ
XdctFWdfD4Im/q7j8jDFKQQoNRNcgpcvUeJaneKGeYyo+HcHAw5zhhQCybcKNoalwB0/Gb+mXu4T
GRQ3reW8ulHk8ssFQuBPoc2k8S1nvB8yOGyBUWe3DSGcFRVF9veL/MM/+a0NaSlqRnULPtffdXeE
aPgrKn6JDESQJhjbX+MlRHmCnF3/hHCAGCaWBmYSKcR30TBy7qKo8WLTXZ7qxTSakvHVpHanXtUi
YJBTlrZb2F4tujbhITME2jogB7mSLgx1ACCuJu1w76lNK1AvTg4jCqRprxjNzb0S8DRAWNndpo6X
mC1uGsB2SoLSsCE7wMcHlXu/CUDGwRO/e6DEmYdC3FzPq3qVEVNoCrh3oyNuR6k+b3lhfFxKYDWC
hpjt83lBk/SDezoaFdm/izQ/PL+xc8N3q2MabtcbL2J98JjSZ0SUdXRXATyBVZ+/mELuVuVi/p+t
k2/VUGSoR+13CoGzmTz13leGeVtyaAS+RXtudWb8cO6vd00TuP2l4an8g6Gx75UxYIigJrc2eccQ
6kOCWMv/cTYcmMKebkJuNcTj/aQcVJrsIX0OFbywokEb6cTenTXnNqmBVLt8q4WxgKta6Qb94AsE
J+e2JTcyHrX8Wa/u7t4cKwEeKpriuKOv2SBKNoW6NOtXk8Z9bfRH0zXCywhmrBrB3ndSqs296hQs
pRHsw9W/TXCiZ+1YSaNoSB3x/vIoVnQMO8yYPEBn34qvmcQvNAzEreSXyPXfW67PS/YMWurAN1eD
My/2tkdlZiENOEQnvxZ5FfYwE2V5o5+iB4191VCt1mkfe0qaHdNIiLpmJkr7KAcTYxeBaSuSU0/o
EDPGhcdCviJs9G0f+tJ3qaGONvZJ6zpHukGbhyF8cbDk/AcdG3T7Ifi0lgEwRyvJBIlNG9joNZdU
nmDEHn9UnOg5R/6mYvf2C+AL7xWbKa+jPGpOyIeWZtY8HtXegZxGNMBiWNnsQwhTaX81NzA8R08u
QS2kEXHvUe369Y0hVyWjZdY477gBXy8vugQqCsn4sE7NyDqMyOg2tRd6Z3252BvjWO8JrJXykiXB
CR/NnnS3vo+hj3TfwdjR2RkdxkObci5Si4OTinFjY1sM49n2bz814uy36Q08oYSzptkNPQlywAxK
eQrapQjBHvPdZOE7BMEQieXn7WfypqNRCQ5xYsUxNlEyb0XeAgEk/Ht24YUcwk5H+lhiNW/c0yuB
OPOlhZpkRDVpC596wmHQ3pHAJWdxV60d/RUYQbdOQN+9wcFPE3vDjc7tidjWcE+bLWTr4GcRYMC4
DMjEO5LgkLrUKoeW3gdVU6bPu3pDh2PcwAPDUKAN2kWd95YfG5JKK5iPMn2M32MDMlqOoaj4mJjN
CAMasIOlIzpZ3hB2WI5Nfj5OSEXs1u+jMGNIzZgCmVlE4C8G28a2ICbMxWwDhfdFVaVKvqe5Xqb6
prrqANLWXChHV5wJqqtXc3ZiaRdtboCelq8swYPXtfYuxiu+iB623e1sOESPFEVgZFZACa41V9uG
mEd/AndT1vVycWT7bgLznCEx7dYDsdw3AwlPmR1/0XqE+zwJr2e+TsuZcqvgLjim1eqeXVKRAtQ2
pHJ17u6shOg3z6Xw704TVADGnMtSZOf8M89af6pTsazDy/CJpa3fqAQJbjl4uriHV7m+zKCweBQR
YoXvsUYejF/9O6/S/IKMG39CAwp/CIaXm1U2/eKdWlFOzb8vDGh0JdhQZfoFMce9S3UvVzOp6qp+
bU2EFP060MQkVoFTnd7ae/1TL1gWrFChpDFRgnqoQIPZxZaiOhSohI29wLemLQan2ObCxmPwDBix
wF0BTegiNgTyCY0D/xjtyLn0uy0bLNFwJvovJ2+jeZVaG5ql3rfnHZrn8DcZrxulCCQhkt8tTfqd
O2SQ9hibT9vdYJ/fPAWMfEzo5oq4s5KdjN+IOyIfjE45zWBvwn1mNy//L5Mjaus5CLdTuzwZDY7i
ec2Pz5kt0Y84BOrAg8cuxe4fdFnQt6xAkXX5hpvJaEFIBfyfQpb4ojgV33R9C/AQwXB+pf13pjaZ
HkOQ9EODYY//9lOvY69PKzGbapQb2azEYT5KpcFV15bfLQR8kHkFFhVK9o3Ut0ZBsH09OBwSdZ7Z
vgsVDj5E8CKzNEYOH/C/Uip07nQorfGqYsXqONyFWL7Mq+ds+VgUwguTMvKBi6VrCkXm8SdkQ0i4
KqXp+I8/81qUtlCKs0QpAeBhKvoixsiNWhK3G6SYZGjlpjPLHaX3EAz61BgsxhjRefqYwtIsRzq9
6ID+lYNMYgZ2p/6AbJqAI5GhSeQcCvZCZhSfqCnX//gyEhnea5B0cauAD0IHGXxY56rUt1/P4yoB
qNkkDAlBzp14IQTRX3nuD/heTd3T4wGebqSTdz9CgnWl0D0ny3Oaq5cprkYT5Z+rV81q2/eZPU0L
QhebLu6pc8bqr9HLXWrHeY+J/TLTif6BG7iehR9jQuP5anCJJMwaQE/UwJfeE3pnRK2RpLEAAiGl
LXbgiaYmyLokeb/HMktBlD37sS6x/mhLguIp7GVaqwY/rZzlP1gJI+H96TTljlXGgqrvo1NEQ71B
Sjy65ffIaauFPbTPH30U/h4pTdGSp/nzmPXWtwXQumybnP1xv7DbzarHgC81w76HBptDBd4vSpwK
DxuKNWR1Fi+sOgBGiKWzO3+J4Hi6h3JNdWBvpCFae531qIhwsxW02fpoJ2G/auLOzpo+0W0Pb3aG
3S3u59EgZ30ErQ73T80yR/bsXVYoiZfep3dPSUr/XBBzm9OT5yJY49iXMm1SmB+Nadtnnd8oyGv4
PsrqwXyBtgRUOjaEmR2i3l3F/Xq0IJY2RIBBN1h/bEbYbmuMYpd07ySHepMb/oCOm606MuUB1hFH
KKijqNZ90IdMK0eWHh429TewUH9byRnr+NBERqY/GOSSsGs4up5pLbcouo7cvTpj97gaB061AlGn
6/JrNL5p8lM7c17vHDqx2+6aY4iQwtIKDIMVr4OH7AOwpd+iHrBcMikYN+Wzdr56UxiG4saiI+bA
GL7HzXnGUUYp2B4pQW5kH0P6cALjtetv5dwByRscMbm4F09swu5xt3EITiUwGnvcaD+YnBA9BtkS
E5bq/BchAlDrB4OoGjRre8oYnw54JmuwhMQLa1knDGw8B5Sq9U1bsNEBO69QvKxCSD8v5Ub4E4So
Q5ojX5pUiqPIY5LyqeVRAV0mo2gGIBqzbyYzVmDI2MKGcp8Q0nERC1j+VpllDJGVlyukCTBQpO7U
yf00VokLPH9oRrU15sS9T5f01ILBb2AdHxxY+qxjvMJ1ZHo0attLAXYcDC9yb21QSNDYAJPdFLiK
Gf8NQXuzOG1ka5fqrWFMHRKKAeEFmRYddoiebZoCMrpmfHiPzwuqzVDLO9GeeVpUw123BWCO8k7T
29USf7/9XwdEMc4gGH35O2FTAz2hxO3dAo9o5f41O437UiI3UexsO+ySelE3Lc2dhmI3E8KUDfiV
8Dh1/P/pstHno0TSZEi8U/LRjZJLxckqTKqFQV98phM7k9ksNN+r9SF7RJNzOAAgcRYy4/dRb8Xs
g2vozZefR/ih1SZnxyM5DUbfu7yfi61jBT5CcwT+r8jJQg7syzt9JYFQbt58OWIbuGDK+wMzPkoM
1pNMf9ZeKRSmkL0TNlTONtMI/ccoELd9TAPIMhvpEIMrZisU0i8dDXTH9HomHk3EaX/GTR6yBa3M
MR/WHyyxeEXC3UV6ia0YTM/BSc0pZJN0PFmTUyCkmGd+d43GQ5NEUlNY6Ig++iRQUzokNMYrT6ss
W5+btj0o+K6N1bh1TRFLCqRunTsx7rkcuPzFqoQ8zWTQQEvXkeY+X39bNBC/cN1KybHaJKYnjB2k
dq/dipMxU8pVJRVcrZbkMXiQ5zVkiq0ItCXrqVtrllBJGloWU2kjn6m2+9onpBKc7QZ/QR3vadDC
WU+ubpX960BxhpkRZJLSQ9X1yS64QWb9LGSu3PtF2d/kDoYzTW4dqMgpYbTXgU0cdHdn968aVmiV
5IHQsTw/FldwbAG3GWP32MUM3U7EmFtUlboLpEfU1gFydlrLyQpyIL9ZDKt0YZCdtDeIJuodzVGv
B5gu62clgGDlgirRT9NLfyJksO9zKKNTSGQ3Wd7CuehiqpeN4UVDUg3QjNCxhC5TG70zZUk8xnY3
eXG+xKgUX+XQOCzSzSKGYc7f2UyaXBFNy5YbEfQnWi880Q69t/ug4lz0Jzoi7nLjiYA4Rym4HCNU
6AHwmzAFlhpTnzyX4Ef8Y8hebiElkj/oyGVZrAPrNBqPnp6H0vfOFsDsUjncbncSWNr0WsiHm75/
YO2KhC0w6ToKfZTmU73y93ixhEusNBL6EYPLcT0MDuPbDCarmE0Rk8+3wpi8P7rpAotZOT1ecyVq
vsC3zPb4HRbqrosOgT0n17TgC4s+FnM6Z6KVLgX1VKkWboZkZNpED1DUmg7FlUhf0qHwP8qbvtZs
Zb635X0tWx8a7EHkDtsjCnjeZxz+KVytH54rxZrSdLKAfnExkz/pjed5yogKuPVLqEv374KmVzbT
UVAT9c1hOKMayIcptAubvg7kbK8k44a0Ob5D88UbDxmXyOBn+h/ZbRn4NwGNyWfyO4RRbfoJ0kTX
TEjX7O/wb1Fv9EujVShz8BctvuBjnAuvS9NRxlDXIiVblUMdw88dfh4yHZOgUptDo5ncpJfbuLWf
ir6ORYlcUL1fMongyzUZBSrWmc8dS75UE5EXYZ1FUbLgkbBCf6Y0ydUI7jKO0JGN8JrqxQAJN3QZ
5K6+ccwH36RuStgs+95oRZ0u1MIIpu5TsBbgQ7PqkMQtvXHtYdUW6j2obB/7hrW+HGwtz2hJ789H
+kK7Ze8rsrcjHwx2TUyfuULdVZE3//O9ZR+i8Bo+wSIdkrTJiJ6AG6pRH2h53768BASWfUWPPXfp
9POvlVdHaTC/SDnfr2TbDd0qecIJtPF83m1afUzwSKO1+1JPHRkgL47qVfwzRv6dzWZ5Btcuct9U
IJwQkMSEXo7VjBSpZCoB0gdHm1JC0CR+DiJNSi5AUANoJMCuZe60fTwCc7LR16WL/9v5E/+wflKD
uFv584aKs00qp09/gIY9WsylazM9omHTOsgce06C6bA6drS9SLg9LT87BQt7j6lJQ3MGqFKSojGm
GMXPiNRNo9Qiu3NG2zRUSuGbucLQRiqBLgldbQWOEtjNKY8JSfQL7ozuZfN4GXZyw0c0GWPiNlno
FoVvv2kxSjuKj6IwQjjOiHhPxvyxN9EfB3U0sdnN+i/z2UXQloMNYR22lawzeesLT9+qfTpJSZTT
JprPfzwo8a+qswIV3B+zjGcJZo9wcgegZeICiQ2JyHCbnF57ONjdXBpSrPsRGE4+9YkZPe9BGDLC
s8UjqSr1/CXeOOqAkq9ZdgHmwWqy0boBx6lyBtNu27qHMhacxrTELhmXUERGtNpcqRHyNPYYo8l+
lEgJ7BGP0NNQQZTBF/5s3h8Pz+d2904t6P40TtGe5oMs/Qd0U5T48D0q7Lxdhin0Cytsu+hn4Cwi
ZIXldse9X89BKVHXTlc4eW9phaa4JThPMHmYeTCl/yl9gpMijBkpWL451DSiXTDA90k+3xi3iQKc
2tFQ5N4IGD8eqFcJeaf4rc/QrNbB7GX5ovsdUEsOG2Jhyn+sRAdM/mA9EU8i+sJeElq+ucP1Rd/1
7mAsDCo01wIUaezjsKeWhUltUeq2W5kofPcaGOVePNt0/mcusRvGry66IadHn/2JZl8/5/dV3eIx
hk+lpr54Th05oztUnC4HMi/PFzVHXPOXMDE7OnVL2kXfVFeczyx04SODmTVp/0w+4BRJM2DNL1bL
OigcW8uGDRHcQJBsB7WCWJWDh/LYfPwyz5iLl4eQfNp3xk7ogLmobG6AGFDq2PMubwNOeJGDoBmD
0Nvh16kGeC4hkoavyyE0ozjLIu4X7tqXSoj5enbAY37bBENCK0YR/I5/vNjfhsM2xuEG3IrQE6D+
pjChi3s6POUTOh2PhZv4epZRsvaNej7xx4gW66WVZGm+ABenn+uKkU2hkTsj4oeLhRf8IcWJTO3C
mIfyxcKDOB0+ZmVuO2ntcKlvY5w8fZXZfZC5VvAY0DAEGiiR9D+R2UrTl6F4grEdoqS5PvFeRAHM
qxKDBclhlrCqsru7EdqOuiethQ6aVddDTjt8J7rOkAhNeh5g54EJpog0aMKAhPXnM2BxFgWfuY6S
lZlGIps4Koz69Eotv2mbmF6cbmWdDiLl0y0ev6nJj5epl190ZOOEokFbp9Cf2ah4KzdKYf7+vyYN
YW/5HZ6frEx6RoM6sA/oMmYa68mKliF+UdNEP/TXi2iF77P7d9lo6lEVAKKSbvP3+IgjU7HESyum
gGaeHld5t0Keg71n7rfzDrT6CdRK4K01NQg7SxjjAxz7GrwLLcan8zqH31Uu0C8PiKwiLhtcvdhL
l0aXYAz1rqBMj5vWvezf+Gc54yK9wd6xm7pCios2mQ9DBFduGkDT/s+Gv3IVJ5pf9W+DqDx7rK61
P+QExj8u5WS07zJ8sLLbJKxpyLmH4+2QalW2DB71sMfeUwTPx9yYG7ykmC8uV5kKR+AaLApQKRhe
dp8pGfNnIzoVx1OKpbdbeTiN33jjcOs7N/u7yTuOqUZ7B1JdJY55m8nM9+f7EHrGWe8+rk/B0Exx
+flkTQ4QUSIiaj6k+e5nDiNMkvK9MoWH+LMrOHmPxGBKXhrfEx8faSMZYhKZ28vNZeoZCMlx+nx0
d4mgA1TXcFKMzX9kkYmTa6KGkTR1BloOdvybUGWFqKTnG6wYQadUF3wz6Fi/GGI0Dl3hxwht3KEg
EqCKxwpePXJeszH9BRnJawnN1wOZrEtPX6EdzTjl17cZxUr4ZjRcq1tvQdkNeCKEEbH/GiO6VQVF
XyzeDWjMCSicpMXV7Vz4JlhSung/DFlq5XdVIOEwdkG/G709rq+h3l6rvZb/XnXuKL+CpfBeX6t6
/GeqKLYahh7VWjQUN5F6Qu4Wlz/tH9K4PtX6GL1WBUnaoJxtmDSnqV0SP5AhzZgEdOxOlQmsckCo
M52Wb6NWxtMNz6q5UPcL6S2D51gLScoP1u5yZQpkskAPqrLU/sEg1u7KmTLuAtk7W3HfqYYnsgQn
5U86pf6Oh++fgdVKqQASHF46/W9u0FnxlZaMNt5+e44lXSgLbGggrw/lYiOULKtGm97xXFZ7r+Gj
Iq6JpCEgEk6Cz5xvyjKHhRzyQ/KS345CawhkFZ7T2V4pSnEEhSSsS5GkEaqNg7G3ZZFPwLzug4w5
xPWgsr9O5OxR1Xq5tkKQmnoTBV3KIcQ7JVF9PL1i+Y6YOdd5E3EPHEM9cAcF5EnjpNZ0/vIqRcu/
CMrx61PoGMXNWm0Vc3PQyXDwcursXV2ywgi4+LESqkP6+vC0hWLr/aUGF3yJRzh1s6gi3QK1LMq2
F1qr69q25pQKUTDxZf7h+cwsM8KkzgqABt3VgKuT07XJp3PV/rGxIY8jf85yd04hgRpqlUhHUr/p
KdyPvWJSwpoSv0igyL+IwtRWBiDATjgFyS++zHfhpXlBa6zfv409VLsdk9abZcHV6Q1e/bm+q+b0
kxdzOCuHpD1R3mqvWSpyg4weTC9apxy/hbgG9aKC3i8umjlgCqQ2qnGAT2E8im5sscHqFbl6ycER
jvqcb+GM/kpdTMJk/WIo1kn2cWLEHlabxYOY3MxVwgIjlo93kdQl4NyBc8u5FtA3DywPWOSvaqu7
QGeAF9fviDRcjMqiilCahH7NsiKSzVsfpAg/MqBCAg+ElBHYU7Cs6P30xkr6XdMG7YdBFh0uVq04
gzalTZEkFItJOBuf4h3JQWafqByST4sCRLhip2zM6FcdpviFeVX3LHKm+4a4wLlRUz/SktT5C/4l
amATbHX7LFzgz1s6Rcc7KCw0vb9a+MQDcqEo8wx5QLd9v/W2yTiE2ZNRdxWNIY6ZMnj/zxNJFxe3
4bV3JvxknNqpcwbLV6M8MjP5Lv45aTMMOE5V+u0/xeXXzcXa7CZ7DvlChGfdbYooq2l7SSCrEOg7
NCZnWhJPXCLFszn7NEZpInyfjmUZkw3p8sjMTUOlZeYbp6qjYPawrl/e+lgATapXJRtZHqOVk0z+
e2MN7SUPiSyJt/rTyzphCiwoOI46Q93rw9BCrPF7XyNOgkyOPDDrWQmMCezG+aadGyqzn5ULgr2s
ME8A1PZsMpEBGZ4/W51kezwOTPM9nVujXjdENiW9Lwj/BPqS/DMAHLgjVLZaBLB3OCxf/xv6IVyi
Nk3S0vI31R6AeubIE7qbxzyR1RbpQhB+k9sE1SUtrEghaLdy9YnpNd30gJbxGblRAByhGxIv29kX
GTW94muRHnzGCTaAUh4Vr+MYpQAyAPvVxFvv32hbJ5VEBdrO2Oke0KswmpLpYHAbSVBFpfFUXNi0
zKjYZGYK/NgWMdfW9ByCUn4qcseZ1cfYJJDkmi7XcBtv56EI2b1xwikGyY+7EaGwbyOR74Y3AaCv
jwEU/9U6qi9XpOcByryi5kEi6on7CtgQBF17BTsobzraP3P5dbjFfbKKL9OpuLX2xnJx9gUB4Tok
a7dGp32S7UB5rYanfHSj5WlHOxozCKbmgViZ1fEtScRl6cPJZPDFrYR7peut9YQrcwKtZIa8dO2a
LUiJzbz5Rvddq/VW8TY2UkY6LvmFBN3FRxNjaTU4RJmX9yqwCYX2WkAAm36vQlVOvxVhAX2QWogo
iFHX4+o7uIMh6EkU0RrQYgL8zd+93f9iSQkcDRmxfpFCReFbM4p+4H2dJkQnNudA7TqLTmJvHxRZ
ibtC1azWGgkrV5qIPo0eDONtlhr3Wq8DYze6/jpyOPDkzrwvVEIV9PN0RkSeiRDSDuwZUbXMGgy9
O33HFdQrfjtwgrkv0kvI4UPL+uJXLD5Cr4AuJ9Kxr3t7455HcR3s4V0b4xfjnmwurMNK6e5vE1vG
dm5qCfEW6shcXcEWJk6++Tf8T7x0Yr6Ywyj8Js0jOIB4+rbOcKYn/rjpbMZty82kFGYxz1kDj41F
zBvFfmy3u77JpsgFbWU5GDeQaX9Jk9ddQCnh8Awlcp6Bu4dPEkX0bv1IC6WzmE2MZ3hvnaOPcz7Y
KkJn3HcKqgau/oTcs2gMkJkPCwRHuiIfMyYC6qRQDPNuRudxkgwP8FoE2PPnXfPuGIhxtnWAIVfZ
h/EwM2AdbQJ/xDKEmu6nkqdJVbHcKbtwpOf5qGKbKIIJyjS3WLhKT4IgH5fum7NpWZ2Eb8fJdAb0
VQByMQwD6kF3Cs0kkJkwYCtwzxSZzkuAiYazieATJiG8WeJlySpYs+UiBCqeS3bSgAGRM2PZji9r
C6U5sR6DLgNxNvIrdID1ZQTqusw5DFEwwXt9sqgB+R2/tmXp4veR7Jm6BHV2M6eouZ9/DqlcAWQU
ZIOXl+w5KkJ4e3SPSoAtorVI/r3nc8DbA5pwdrRKt4DLnkIrRZJ+/uuL3OuSaFL79IrJywb0NmOq
FwbWUhjaMDyIutEjH6CiAiD80OpBRGuV3bAtFBwXZAZQXW5D5PzGcKmW1cdNOnvkI9PXtfb7Ybr0
4zP0lj4CrtzY8oQC1xEOrO8pnZs03H7xi80mhR+cC9npiJvT1Y5v+u+ZHKuRAVFEfv4p3CfJdA71
Z4Kfuk+j56X4iYWTydgZgxqw2qB4mo9TMFn23cPh7CHc34J4bHKAUsXnSncOgu/P8gwFaWwQ1YEr
r+GW5OTvP7Dq7eHYblpUUGg0JeWVAbXLP6BViQ6P5twYBy0JGrim/bV4k1oeUth4gRMNBe5lCcXX
jVvg8CaRYUtkppqlWl7KUenqg4rTGTXKSZElkM25g8Kxc5yXNiNSvxfSeQOCTtwgCoi6BBjvuD52
CUyh3wJRSAM+lwi40+gGpBahcF5xEZ8R6B9GWp0TyBweyhOGKD0dNm9bbOWVCUxc37lbvMXCMLZv
nvWhB5V2e63s581BFYJlq7NZP9IVHWEI4Jhou82pO/hH6j5AnHXoLsxV59kjfzpa7/PfSnDzXOd0
QXbCASxFYACZpIgf6MhfGr/HcKaLQm/qSFaF5CUIXgdn1PIOEEgz0aHGhbeSTx36l21DXK3p53v7
Q1lgBUiM+GvZ8sCpTfrYJarWKe8GbiSEInCvg01FRsdrAtJAxtUm2FvQlXJzpwcqUK80FOHZxsLI
UCkfBkINE4APdj0nxU/VQEm4GU7U/AdyzIapreR/lTuKt4q6pWq/zmH9mfcWvaosgOgbUaKxFY5E
t5sx/4mTndXjDk9Jxg1zmJptkrN902FfYSNXVAHuFieZDuL4N5+RNwF5kyFrkythIJslep0Mfm/B
EPBALUVEiSgZQcjJEUwspPhBlEYjedtzV5/to/Vr8asmbU3AtDzvf+n6pDx1rP8ViamebOuFezNZ
DrhaHUDBST0GptXvJh+sK0KnkQp1mUS8zHRckoQ7LX4fGXJmm2KvZb7/4W4d8qeAwYiRX3paQCYE
2ybKpH3y1tWLYX/V2RXTs/6WzAGAkHHaC+8AADovSIXWKkEPU7pUIoEsNhxhpIW8xUzqAlAZBLGw
73lDDWt4frPq+909Vwf/GHKb+Myq+r4ht7LZzbtN4IHrgdBnE+QRN9YARCeqzQACLCKeihKemmTY
hlovUtMKqB3mGzeqnSc5bQYPbU5W0hyAx2Sf73o4GmmKt+0bfAp8A3FZ93AV1eQh8Q/muZy5LOfT
hXWnzY/jjqccc7HNzO4aoVqlYo3F54sg2bt1/orbR/JEEvcw4AMVOwiKnWON2fFu4drPnv/oZiOG
vXD0S8pj5jLd6Zh14o2vHELN/8GA3nOe7Vfvv0TMT4mPyDCbndeSeP4TC2JoslCY9gE+QAm204KS
RRE7Xq8kpmH1viAtDw/6ZqJM3bvPUWBEfwxeGqqv6Qr4hI00WAHZaBNhWoxwC7GfDSlBeQNu+YRk
KhbtlwJ37+nNL1QOypoIXeSIUoertypgvNsYI+UYQLVP4bbFy4fgJb8QMRhPMiFwiUqWUIxdhcrK
wDbvXepwIjz8FpxB85N5ltV7tNleqfcyKV3m6ShmD9YPYE7KU2zh/EfvslS6s+HSQIhugzvvL/K3
sAQMaYEyuIA/VpzzvzfSImuD8yCOlaOkn0n4DmGRMiBDS56YRo13wVHxhQ1EA+3W19ZmksSdEmf0
1lZ1nRFr3nytnHWFn07wyI5nByMggsuP8mnZAr8H650h/y2TCMIfF5+hT+UgRMggufL8AsxPC+zb
NFPWZ3nxXK7xwAuIQwjkclBrcFxt3HMNpAojTe2oPpfFKNJtZFUkfIo8A+zrSusVknCpZeLTAN3X
5WZXkEL7pytGnHGGSrRXzL0IieO1549nBcAN3MF7EY35gtD9deaiiRdtQWjNFEYs13/Sk+GMIboy
wDJVBcj4LyAbWQ5jjWSNi0Owc93zH+KTjGlxJmcwAJ/dveoUBVZTc2EC6aRl907sm+Bn9HHLfDYR
JcTBC2FuTUbPxs81UVzJNPBUzFTDF6FjdY4wQDxpHU4yYkg49zXlHPGilwtGVG4X3aT2ajURL4Ka
+5y1cKQkQ3dT55PTDYWVZY6VsaoKv/+sM8+bRM2pI8c4YECCX6GpDQ/yeJDlq0Gl5Ojp5H/JXudY
j5fShWpzVIX84y9FErfTM3pWforTKUwBUfZqxSMnrCS07Ak66hgAUCt8UJOD13zxh93xyDN842VV
PLIkP/huABiuFXm5lvSwpPkCN+aaOzG+nBBA1+9gST0EO/MliNhEVTbZo9O6PkBKP/gRVIy2OwT8
LdDmrl0wpBf2/AlqgFruqSFhom9xeQEMzRZuDGX9Z2ME6eNTN2MpAc9c6gGFToIm9Ig3ZWamO0oj
lXQJaVIMyNGNR0PXYOa0qjWuTWClsEEjxUUi1+g5zR8ETt527FqFf5u+CvcJ7Hhh54eOSTr5xQKQ
4OSDkVKhuq3/HN6wVqaXAkZVBbXEkb3XuHkXc6RqJofZ+Q1HDHYmOmzSURVdiJrHOs9+FnI1reGx
NctC4CP2idBGfs2kavEdqi5ay2m7M0Tv6tQeug921AuaUVhYyAc8UYa4qR9ERK0JmhKquPQ+eYdD
uyU3V33cnNv+qK3j2TvusfO4l8xTbqygLQRwZ/yf2+cW9JZkhm/xpNrdoCDDvvyOo3y98LFoWG2j
YkGsDT5zqPbMyybCnS6isNAK1UhgSdq0/Y67sdvLmYv/kEHy9I7pV/wwv5Os92RieqQCfBgZn02V
9ZhdiM1a0aAgxBWL3zz2asKYYss5mNQvCSh6eUJkG1bJax2wh6pUyAGfsNPgc3uXKMCFa5g/1bcq
XLRn23m5bkKjpx1wZsRgToI5+vOxY9R+Cbxxugg8iJV9LoXHul0vxop+rgeeuNUWtxYljNstSoVI
jha5HsjHMMiVRIHzNWGaqyFCACH7sZfrvSR4oCG/RaKugD3ViD11mrS3jcK/L1enHeLa2597Prj0
8KM0p+TAds0wPtZNHS+Qar/Avreb+qYshopMJEN4qdq+90qAkDlvCvYSxiVZXZEddylSGZgJmuks
JZoDwwjmftSTPDT7rHg3chCZRNWEAQVCPqzCHqh03OgQFBRwSB4/MfX/Qourd9vVfkuN8c+J6bL8
Z4/6Jd/meOYsKTJ6SpKDBNQkuXJBwF+kcyP0kDtZQkHgEMVTVJoj8Q2COGN9psU6WcL6DjYqgu1j
ifpDavEScdgKlWEAvihZtA/T7ji9zxwYtdcgN8x1RppHBDgWlnBfAqdetatPOi6D0qEvVWX4DDwg
d+wogONzMzNb8qgkk4P6dHudY7yXjBEAhXBVfZbYgT1XiaP6gqdEGfEJWTAkkWNPkbPFBQ5KWx1W
ze+LBcmqP8F5Foj76I5rx9QaExVS0SOHPiaymZp4vulpLXof49bqna1ON+Gk2VhQvADpWqBjvnOR
BeL+ude+dy4/UiJuyP5cSWfYflSE0i7He4WDaBq7xKuExRBbcMwEaLHHQLb9WpTAo+CAKHiw8pLt
Upv+eUlBartmL+wcihrYX8ADQYJejcIcwZW7hSfNzDOxrjhEiL26oIY5aLIo4pNvzoo+LX0Jt44n
9wX8NIR733fgaCGbrXXfpztPxXCuHbUkTQKwi4Xq8SeKweyIS6Jw7EXKi9KLPP/oe1OHmT2iwNKu
bgeaY1lUkNoWjZHzFi9cYxhXBW/eJR1sIxkfGLSns6hUqvEhIla9+lk9kbIQbHPBkVfgP42b3KAU
zxNk0SpO7gSUDWgUcMFw8yfNJlC9nQOh9wrBMxnhw5slsCenysr1yuBjQ3SJXtOn5VRcBN6WOj6d
qMZhQlce+7+LNEchE+W8TqoRnZardL3DVdRZ2A8/qep310TCn9oQKcUboJM4RkP8C87Z9/B0KEZ6
RBtDRm6Og74a/sNbr19CriTB9M52XywAeQzm4vw8MFFeUoTnomlYUqVh20+wfsHQckf7cmybyOWv
1wkmwgT4AafKF/OttSn3T0qjElSs9xgTzUApn9kjaXFCtK1ChX9X/E0dZfOclsuQV5t7kBDe61Tc
yMLShE7NUpVYnGZokr9UT9Zu7tnlWvcmsj5bYKSZ24PP3S3mSKG7MNFwDJOyACMyMMCavpwmb7R+
xWBTbLRqpEjElQUsFcAnV6TXdfXH8XxRJDCJsusxHKlpdg7/UPt+M/muOJAPANPdEzITkotAxQti
f2sSQ+lyUXQawTqMh6GSrO+ScIgHwwvZkk86bl3Qa5QtwZLpomNvdkUliHaVDorZcBtVY94NurVG
pVj5JoTTUMpyodsLAhSsQZnjmt2eFyYhagonTyAwKOBrmOZogYtvj+zpsAByJ0K6xuZ7R9GdpACn
SjasnecDfa3kMjUZjqJd8zKjuBc0KE8xEfGrOKRozOFELU8TTE42sAhSIm6RokpRGHXRi7qDnwEu
1kWuY2Db5I9NulXO6C2hLRyJQMOXSHfiPTNgetZOpRPTbvvrnmOWJSppzemvLEDk9a7ghAdrLWug
Wz6EJRnsC/DTfO5KzPFtXcwS1dgO8IblprGPQ+wYNWok9n0aaw6Ic/RLjwk6LhO2+lL5WTQAf938
HmEKQBfOB75QCFM1BwD7bptsgbb2ssbuUQGdUkUUzsd1kEuDpXnqABHGWhGKgv8lXWPTAgHxBez6
uCllCw1B0pMdYloAIXUjMyGJB45kazq9JtYSYeL+fKHJ+B/SFc7GjYyCe33q50wYDZWT5cHw7oTS
yx+tv1j2YYMr8SGZUMXBfXQnG8lVLwz2A4LQeaXQgrCQ3pjLjFphzjrpJ6zmw9ArCYRPd0x0OcWR
OtUZBe5O8Ydk9LlzBbynRHHHgKatXNlSLPgEQEYNglzr8FXLVDaVcox0Btib4j8qJMu4GALr7o0h
+hADK5aRJWJunDT4OAVUYF1URBtAZR22KjxFajqJESdZO6NLAu6h7V73UDzLgLVhjEUPI/D2vcBt
T4urGCbgibGVhTD5hnUOOdufdpgIAwiOQh1D18q/E9sTHoCPIx8Y6UhLu5R4ygZNj8HofC62E2Lg
g/AMJNksSIq65JnwiLgz9t5uj74gk+yrCHffFYMV5rCQUjVtVhzU6N6Sycx8kdEFWXEblmU+11Pt
FAIfesIv2+pHNSOUVANnnt7oh5vL8sfoPUol0M5n76J0v7TW815JMOccU4iGdAfhCgwdZtxRo3lk
m6w7GdB/wFyMB8BZL+aA6/HcleaamCCtiMa2TLpPEPwvMcj6zP+PmK+EnFfYa9Lh8DqtmH0ofnor
BMUpZUN3ABXREwwAeB+/pd2iQccCpqJsvIjhCb8lsHI2t9aQEAjwRVklzJI5pi3y+YEg7cOZoVv/
ko7QcREPjOUE8Va2d6JnMHUAnbEQUw5w0Oy10OrbJOeYWmJFMIkXWGtz4FGF87WAFl5hOcfCTm5w
cvXQe+W1+qFhEB6KANffQYX0pWxyCe+q8bh/d4XZGIBbhrwt7p2/7RlCeoICb7td8jw2xj7aXmRN
+hVJqRrE1QY0BkibB1b/lI2wN1MgkweImtwCpHiE2b7QNTm/xqfi/rzAaGpzhGT7tbhzi/FQZUTr
LXzP8E4l/bd6vAXt79bfXqIYzFNYBYak2hCom2QKedwzGgymLe12xg2fDpsr+nerpn6XExxF0YV4
Zdtv/gyFWJYVYvjyfHXo0uuuL0kfq9My7YReK9Bxa3Yqz3EAe0E/FdaWDaXBNg3Ai/MLDsPVLfxR
CbtdhWvNNjQpY1XpjECY2y4TrFxAJ0o9XvFQtH9gj39g3BdiSgCPg5d5SBgO8S7ovg08dpWPuxon
64285iMK9ZcHuIxDj59ltLOz0pj4xVlVMIh2xVJSobbI5hQUaw1qZjLIR0cboohIi6aVkvOeGzGX
nauqHgaZkj0KxxHagVamhwaTFiAIi1lmyzxkkYtLZQuRF5ULxG6Ik39N7LR955ECz8K2G1/lqyyY
AykADCpUWmbk2ZqrK1xDdJfZGrPTid/ZM5mdf+kLWVJtt1RMUbvlMr0ybxxOoDoi680eFRjGnjKW
p1K48VNcT9wsWr2lnD2ZbdkgF5F08zRkFbhSnXTNSJllXYukz1lwRrG8klo+66cORV91qozaR3iZ
QkJxHHBI3eJOCAxBxUizIMFxXE+yMNFoz/5WYsszjzUj/IIdLgLnMcHaC7/mCD4x2/9OFpw2i16E
5aTtcEshtVBowwxpYfBbmmjQiE7xLSVmM1tTytxsgsOJ3xz+5smokX3hzU1Ht/TuZRcozGeec0G7
xFZTfDp6vQLQCfTmuDSEgPjTnSXKQiSEMz+09++JLsQ/Mum9h5g0EEyOjQ5igy3e4dq2ZE7jCvxF
EVGO4X6iJp5AtQVbLo4iHVLimM5ky4QcNI3KMdOkjpD15COqHJVkABaFI0s2LO9ktwjlnA9tkBmi
AkaguVZWT/QkVJLp97pB5W6/TAXwiQuCDe2I64q9zW7A0OWco4+B3peT85WqpWXq02ovOlgEn8jS
8afpjvCdYrAVH8KM9C6YFiiiK3a7HTeiNFSXzty0Mv+5cr9zfEfnig4wK2/VJrIDArru45z2X45V
dBxHI/1/GA0qIA1a+GRWYHVCNYOAtHEgXOglhOpEHN9/AC/Nrk7U9K8zRzGA6dJejM0a2N71HUQ1
wLcNFQUEQkrIXp6MelV0rlWZ0LzzFGECjzEt8Ppi2aqciM1ve7lMOFHa1CVWhChkQh7EcqjDkkhV
TXMJkYFtRSJfTQ8PZ8B+/E3eG0z3v3zZo4o+YNuRbTa7H50XHFWHg+Tt3zks48AOsC1CwVxZLv8q
gntpyJAMxYPfxy/KIYxraAInicpC8ZNpdamlpR32gOJFQKacucjYNtdHxANwVMWycapKNNWlKDm5
BmwiZVjnn2YC4SGbJ2AnDg7j8mqPGIOQe9ujOJT1yXnvbnRtvfHIEv54v4L48t12Dhun5L/F96UO
v2eM67SS56tlvLNiYNmGxMPoDd0X+aU9SEPNf5IIt4VzOEfEPqKQkQ65irx+oj763Z1Kw2XNwiV2
M00xGSz/uxv83lVUkJkbUo/GsTk5/ykhzsKEHYZSQKdrx3mAXE13kG2nI5HuGI6UBq+SZDOHfBbw
NsUElFbODafVFZdWmxHbyZ9MwqG2KYUUoorc02pbcSSa0Pw1WPM8DQeVfIji17kCVPXCM76/PGLl
EeP6oje1NtQDQouX+GmMD5OJ+zbA3PGvTDTQObwwA+OzEnS9eZnzii/qlqrDH4CKA458cttNNQDY
um6JYYYuVju2eqx0IPUE9zHg3w06jcGvli2BByuZlG6nFXTJm4OUFJXKrLsCO6wPxFKhhottGo7Q
gP5JZFHnuVGX6iV16U4ISy7424PPnBMbcZpI5pHAUm3cDbnFj+q0XddFwndhABWBnuNQktr3kDzm
OrFlSaBVW4E4nzapV9o/GatlwheVmtWvSLfD3zhqbnUJ7urNLOCALfWxYqGWU76PGhsQkp/gm/P4
uEdcYTvspQ+02/7RQy1mlEiLwFP/4ZOxvpTbHxMQk+IP/Razk+dKD82Ufp1YVFaTsIg9GM8Q2oW1
fPE5dnbi6qEB82GcE4nOcAqGcZTM8AoQxdEz5BU+ualu0nM+bUhYcnxP/vPAuP+KN/BPAwHFZVyN
233iL5rCeF8hSOp5RXwhvk1vPKKFMZVrJ7dHrXGcZBrIycu7yY6K+AL0DeBZZPUW0WXQxRA/x7Uu
b7951bmVOFiNsnGnILbdRoxOtSvVUT8ESRjnoXRcQ20iKurLqwW4L+ApIXg4Sb+2RFp2MpvDEG1l
KnvQNaUfsG5O2IXLE1FD5KmlILRjTv3u3E9GVR0mhu/Rs3hmvkr2PRVjAM0Ic3pBocYg432UR6Pt
hh8WJ/4QabUvLsw/WVBHQDviVArIeAqu3phbCue4kF3cjTZjFHo+SyKLhtnUhHjI+mJ/H93Ipa0w
T/UFE4rPQETfXJzkK1PvHh2NGKY8ksssaeXYyKTlFQ/dOiW4+AQR/tKhSDXzxoCCCrt9fZOAu+8T
QOWrzCVTho92GtlU5nMX4wenvcLGUqEKx7Xobk1oDvVOkU2IGb0GaOF56ULjsF+LPpe886Zk4waN
FhaBRMeqYQQDGz4yW+twClgdx8tUNf1GghaKukVjcVyaD1XgxXze/pfGjZ2FSYyRP7JQMRaPpEZE
rL5fvgDDk+HstOdCM9FzHbjI5Qvgos0zMbdSGLB5CsvhTNGCNQyE6gJ1qfxcuRGz/bYTk9OVRJBR
OJ4PWm4blfwTUNPfvqpGFUAra2iK8TGnKVa1x9qAChMMiKGxgnkj4nHg+YDmx3gnA1Fcwg8MuJF2
mWlbfxTD0ngni8yd04afNVuv9MVwgydG+HlyfYg6of/l81cabzQ9wfXWpvfUn02nWrZPyZcmXxKY
OC3UtQsx14V6wjyv7ifijvNPPLTp68OiyyE0R/YYIkPmwYYbzUla/L1wq4C5qTAzm5cwhxgfWlpK
DBZcpXRZIao6uzBwRPxPEBsB5OJFes79m8+BkU31/ECH1bMldGtH3KltWuBkC4hnlcz8e5j2GsvU
7S32WGUtbsYZ3VfEv/a/pSo/GdKdgx9M7M3ursmTr9VK0tkrvQ+6qCR8IpMcsPjntgFpi64MIE0g
sdYYOLJYLuaEm7Adrrq1pkVvctK1qegKCZqIZc+4SBYsa7NkIPU90TijBl7UGrHNcvZdO9rCFdce
a+tJS/0fR2zX006DujM+nWKILhKdi5mtTUOOmxxCcMUWowmNh1cJDggdNDhM8dR+xez9Pz1BbyPF
hdTPUqbNLM8/eZi3PG8jQPSzM62P6VM9bcTjfDb4ZAe9cNyMYiFJEQNcUHveneYGG/EnTpyFcPk6
hRjtpXzbksaPxcD7NsRL2IpQjl1oIve/7wUwrehBkpqt7Iw140YyNeINKpiH9JyXvenWiHQem+RA
NhXeY4MIYHa9p59ldGYH+VOvqaNAPI0eI7T4cuIrnoJ7YnMD6ZnF92qAbTnzIcdNtsmz5/FspUeL
Y+e+BQfghto07+OLC57vq9GaV3p7B5/rSaImkWWi5feLqWBGpMw78ko3ncDRIbPetK63zx7p/+zy
iff2riAFDTadEfjzmOUMAHwrkNvSnODrnPpdjpavR02Xl9OGZRFkBZSXAW2BDVsgnH1c++ZuXGvQ
n28f6qGySe1PfCStJeUAo63laa1ghvLWFcz0hr2bImzbBKaV9C5cmYOPjp3HbugQakKBfkix612Q
oqAqIKhz+oCDBk+nRkS1JRdKRFfXnr8m2yVRbw9h1nJ1MVcaGuyfjWVRpBjQGmqJOD56sJclA9/o
+d47nWJHCYLX8faXx3OI3HYFb32wm4JSr7uk+tJ8Mv9FjGbMww4Hyy91dWi/WYdLCwtiWKoiN/+k
A/jEjg+KXgPmhLwKLnskbc+CLf/xj6xjGKeEPF+mQwpZsUcLq2AYI7IEvwJrKZm0oYGweyA/Q2m9
n5SNEgCHKbsljIn8lH3YfYVcLFAmEiBZnBlrDDeLaIiod0iKS92e9iig0EUMvIBLBEtICrE0SUyY
folIdDUCl7dqyvc4i1gJwBkhR1GhE6WqZba3SLCY+/U6pmvW6Ire3ossCeCcj4VdfJGqzHQR+n9x
87fvXlD6QohY6jUb+xGXXSAe1SvQz7PVt0FmeNxf93k0gMFoTvx1VR8NVa0EothVST+fxWGkU2zI
VAC/EBduM75SoJAzcxf641YklezWmvrOX7LJwv3rcr7+l+3FOhHhggIZOi7CisffoYWmG9D20ogr
3FGp6ZEychM6PDim4JX7uTgLWw9hYBAkYaY9wv1KP9vsY8FEnYT9/yJCnzTULi4oDZRyTBj8D9sQ
RCvzAJcA0ZQNXyN63j2F391Cmlo0T27AxG8V5CNlgLbY8GWhtB1jJFJ9HJSGu1XfZ3Z/7sJT/dYr
KvKFGGiDYNdFDRMW62BDPIIJsPFjHmZ4ixaWePhxuA0BMpkHUqey7cFOov5xQtfXh+iiqVxJrHJd
LWk7KmyGN59C0XJygcXVtewwAdNKtDg3XKYUlyTZT2aCNLdQDlItPsbF2kFccdcfAYoCRN/crVam
gTe86nt0mAKH4pMwT4FuUOfwb5J94ZG/YIkosgC/gsn6uY1VrdTHE8Y2kZWkXYYAFJ2h75fRm82d
GFqKHGRdN01Rok2BxZg+lPbeAVMwsiGLnToBq9j0aMgiYVgguuNTYzEz6JnMhpll4KVg8rtkGHk6
Dd8xPZMVMGrIT5O6uDLgBHG0Owg1lrk6PaNVlSFaODdxa0x0VHbKXWMzMGH+BOSV/yyE9UgJfAqP
icOIkkoIYCubb1BfhV1kmWZ6e2a4YYuEnnX+z1/B1smkPnn6Ogcbeb8wr05fNdIkRFy4Qga8qewr
bYOu+NDb2aJ6GY/d0XnIaLfj993dRfS3b0L/lm7njGu1yGRpnM7UAoLRSRiFdscUyZm7Yxa1SgqO
CORzF0O7tCDtJpVRMgK2/yVk4fTT9fbSOZxg2cWlx4vUTRkQGKLbf22PBWoctiCvvJdNA5st2+sn
KTOrdyIu8q97oRCgsYrX5+G25UYwHhxFasgCIUwJ9JeKJXd1I348lhv+3Xj9/IfFZfrVs4kHL6My
OGl4LJWSSorVYhnFk1Xs+HdmYetTnxQDAPr9xbotf/R+bTWAO4d5GUFSxRFTKKtbiOtw2dZgyI0/
DGbO9g2vwNgC4R4IS61Ozhtg5xo0zhWGyrr7yuNH6oZeBVrWD9QNRWI/gk5sUwHIES1MDJxINsV/
pJ03oaAZCM96CZVHaFB+pccntNvPg92T3/jgnvwYfZrZAuC+WWvLZNBNIEchm8fuKs2cQCK9MpP/
8Vsi5dV55KShD73Agoo3RuqGn9/Ca2WVQN3MBkJYIL8KTDpyZ2mpF6+x5t01Y6S0TZW4gwBWsxaW
JW/5XEXWdpCK4ZiGeOsyh63EHxs2Fv/nUwc2GoYsWOWrsAjauBGNmTR7hTA8PoEUljyOHGYVrDpl
z2VcP8AzjNcyFIVBlZTbzxjI5bV5B3m3qh8ZHM4NKv1FMZWDLbqiWvx7bI4qapu/F5FrN6vcPIrg
G/Tx+/9oPtYY7fWpCIXzTNaWkDkRdzTcuCs/LHXnhANr1TIRALLd5XYHp5eUTffLd6FNGkXcYM3X
qbYc621hCh0eX78TH107gIn1kTiBCb8bYhCakLSTcAHN93/An+3dY1HNFVKA+aatphrLB3blZKlc
miS2Kz/pswHv/Vnk0SnSnX6CwvmklpaoZw9dKKdhqy6m3LCQ23Xw5bygnz/cF4zcQMnq9nf1k93a
T4m+AqIiVzbgy9XTJ15r+2mvsXauHFWIvnrgkyLcsBL6JkRxvwH69ZWMni1b0PRgP+EgYHOtSxeM
GHHORkL9ZpBmcuyTb8HxKtmHPhtYkwWV5xRVasOnyh1P3qNX68ggCqDJpXrGJM0F8Ln3GkyV9YQ7
xwONc7dQTGyJ3C7PsfNkKGSilLffCZ27Ihe1zgy//NfsUuKBLtvXqZriDzcIA2P+aOQyooljIvFe
ZVfV7PKVUHyrAM83CxO0S3Ix6lSthQx2PbwXaUGpO9TB0Ga9WsTSVueO2eAs3jBJ9XidRR/n5MeQ
KKjxsGGQHmAII8ExvHdSJxZ96zqqA25gRYBt9O4VAQcmwEEHrfBFwmW4aBTZryDIqM+Cgm/bXpc1
2QeO+UTdv2/SJ2azoFgNxeEHyGI+2ak0joklhV2QLNuExrH08Vr4aIg/+yf+znsMidTqv8ySzD8q
aipmBXHwkW8pmtyb5lakMHf/h/dkwnvCHHOqDgDFe1RpWfnuDLge6+ldYjafRO+rfkb6qPzFZv4g
Uvc9Bp2+mW1oNfzGmvPDcOZjZzDzQ/OmqkrsBD4C38JtqZI+wxK/QuuIxrnORNt8UJOHunjbd69o
NQ5dBg7B3YPS5LBbPgFT/gGhF8VKxddkEiEdtYsnNnutKaDqV7k9J6lYi4C8TWbKFUGXqbTcWXnz
psxBKNNcxdIB1qGt4sjtp1IdWDEsR2fF//nAqXPVB3kyYiqEoybnE44bPOIq/qe0N5GlMaLg1m1u
1WDWXS1GvTa0MoYEys6o51YaHM/GGI5F35MKFbKa8Ewkb4fasEFBz9pACfPL1HpQWRBuGOl0i1cP
5YSPyNLt8am33uPya5dxKzQE16fZgNWbcsz3bJPS5Ch5yg62tBmtZyyO1p1h65YToPJ9rs8+BnUS
vf7doteA6w5A/gi7k5TJXfFYH8MNjmC6HBH8Ztd+vJ3FFdvR9XhPeJ/qidvLKUB5ue1pB7CdPBMN
gIb/n8ikspQas3X+mUv5WKb6vutTZUKAbMxyYyqFlJZIWo9xyI0DkSbA8p4zhhO+OCmCKvm9+6K7
u/uO3uImyuO9mwyXJL30qSQnJp5kx6NT0PoBlCUxuHs99d3bT0AvEI0vBdzbQWTXWQ63xrBrmosV
1O04IOTTVyD7cSq8aCDfFjjdJq5UNwdm1NewsBWf0EMb4J4+YTFpSdX++MBjv0Slf+vGDHVYSaWp
Ov0zf+Ep5dwrH6yC07VJY7u2nBh894OozxAj7wgYr7c87H0M6450+ykrxEFRzMk7Cb7l8+4HwZGR
yFNyY9+tu81Q4fOzEQ1IsBcNPfRy3QVhT2mYAYfGW9+M3GTv8Q71DlBn7Oh8smQiOmy1e2rOtIwP
7qj9Iuzz2Leij706u9xaUrFqS48ryf+w4b7NDJOwGU8A3LITq7ievyx7FHbdpVxRtKnK6BAeavWJ
xd7gkHmyPRiFPJowLcTGKLkS2qRLv+Bk0Iu+CH1QCjtJbBOa8OD+/dNDY0nBhxy9RynkX3w36riS
sd9gLmNYcPAuDup7CaUMF6/XMRxpFTiLv8jOs/TbpukycrY0D5ST4L6MMF2bsjUgKrVYlk3Db3uQ
8MfoPkmfZzo+tHI88oxY88ALhF8atXm9OkV+QGlNb1K8svAxxslay7uv2g27XZRHz7iYLoJkatfI
1MwOx0dUhC/5wPWnREyCu55/Ahz3dJYkS+AeL7AzAiOyBighig3s8oFVWqBTPQYkxG8cKqyGZr4C
P/AwV3ooWfKe1MgtoqKH9peeeSAN991g7vRmxtbgLk4J2aZneZxSJbBwWlou2S03RYbZTEAdymkZ
XzAZH9aiuEmJ5SzlXCzWSFRYmHBcJ46S53cpTTIwb13fbKG5uE85ajQ59Zs97UsTB8IQC8prZKIS
FYJPv9nyWqdLMU2T4okmel4dMALxvubHfvhTttQ9tRieF/+FsdxZwxaqOc2pHNXABBJ9Iks548ID
eRB3bDOYWM0cI4c0qeBYgnmbXynI8Plnff+igOasUzvD3l9iJ6DyeY1fesFsE4neV/+G+neTCEMP
iL57OO7YtpSnYUTp6QbLQb3tjXtEYddvh6NyeI+r4OItSXe1MY3aYbcE5AYApKEpMr+lGA/xZplz
f7pQ/Q72yzYUTZDtBc5iqbcuov6DIiIOKa7pWyXpNQwKW6WoilFFYyXIKHbLI8IG0u5iotcp0kNF
dMFPSx58LCZliYKcOpoVd78jFaeM6hqYIAEl4PjlPpXVcnIchwWDlydnPQ4VnSgnKuunRU9qTU0X
vfJOmXW2nQNpu2ay0uZAxMj1t/B1+iPeV+TBZV2Qs8RFrJhUM1qsXy9yi8Qhj2a+6FJwhK8tHfV2
WI35v1nlaJZ26hN9IsSIGThV+PIxgQAPXbVjX9YTcnx3nGqPrKy9/iDr5ubl98vghTeRdMgU3RIt
8hfA+HmmmPfOzy4zPYGr4EeHuUN8k9Fl7MLxB+4P9IOE+ZIV1DOS6M5GzyQ7+XCu0vRv6HRp6UoX
al0CX4G2x4dq7hv03ifH/qARAvuKiaeOsamQbdQxFp5LwxUwsfiAkzdX9nmpdWFzEZKmcXNuZM3I
soEjGQ+1v18IZSrw6zJuPzPfxiynHTCiYfhL5IfLDH3dpR/DhAhbd6ws3vCmvafsVPhOXaRG6Pfw
O/I51SQGGSDp0pMNXnIIV7qRcmExcGVVHWl4UI8v6FqjZRK6fTXLwZLKX+bu1IW+Aw+i+kA9pUVN
2zEncdAtFxztjhaCiGDt857iEvjBQR52O6h9lB+uK4DCQMCDStY7SIA9TSzzX3bST6RuOowm1pUO
PazWUEsEGeLbLD++th3UEnFRQaYvh96rYcWmTPDw8dBi9ATT0Xeq8mFrkRM+G7OGPz3qwoOBCqb+
AEvA7iYxH0KpdHV7JTykRPmC7UODDGmHGu2ytcGQGPrB2+/yWWhlJjhty2tFJVWeK3kWoos6Dsso
ZsPqkwNPldiqLu+GxWigi47FKXWY1Id3ANAKkABdcy/I3qd1HTGZ+Mi1B3BthYRh95lA900WrUZx
aINF2fwGo/8vCAK2lacy89EDZpBfhGxg0W/ygrY7OR/o9ym+qRozXk9zKbZLVhJlO7CKWOASfsO1
H7b6ZHg5ReoLyYKJLo63UzCZAFOH1q2HRMG/IV35wBDXQ16Hopg7mfxNNDuKz1syIWW2LonigYYW
MgEt0iTI/iBubhaj8IT6APS/tXk9j9Hbk64j9oQNwT9PdRuSPLthemBnuZhz0BeNQkld7KuSDb3P
1kZ8Jt+cP49SSTwA/Ev7EznAOrHiw9w8NUGbExLnufcQzKVuo0Ftam0PLPZ0qG3Jil/nojFr7sDN
5hE9YTMsom9zjUGwEeNxYSv1h1eDK2kTQnv+xZPI1FQTWtk2UrAYJUVO3rIKhsBBbDK81MfXJV4r
trNglljIqUdGtNwUkQxqPLnigxHx9x7y1fdlH7H3CBlTyE/qTkTD9hrI8fLsMdv3fDA84w53LJ8C
tzogxj3UfnOJ4Jsa38yqMqd2QxYPsTrH2ef6TJ0FFMrRTF+e/wHdODGjRyVnZaRm9gl12zhckUQ5
u3Hk/68/GO/FvflJgK0UPtUhYWbVDOvo7BhyguG0NVLlYSUXnSz8tH8N1+cc1s80rBA6U9/XZGkW
vaaYBlKh4AH6ZwqGnQdipRUFTzUaTNunr7/pce8vLtMrG7IyaDaqDxM+Z18SPf5Ys+R/T0ntgyJ7
X1n8hWNt2+Rlidj777Wt/A/Wzgcj1MmZz3Ata66aGFK7RAOCKu8ghu+3V9K5ZWxXEm0CSV5+hxdc
MoY3t9PU6LR2FqQdLZWfFI0f3zoO0hq0w4c9vQ5f/1YP1pbEF8L0JeQ9wVoNbzbvbqgYMbaXd3Ro
fpViET4JxJMXPTCaPl9medZG9IuXRQ6QBAbJc6egBw8uYWyvqZ7MkC3e4IvPfUwB/B2XyuHqQc/w
qxDhrq2M7Ig1/z1ARanWq7srQJc6ckUVfuH23hpQjmcTT92bauYodkGDJE7oQyuLADrGIXt5PiOx
MB2IDryjkvQvz9f4Qsg9wtIOSr0/MXdnopEknpFYWo2AxmstJgONGz0Gz6zgO3Dkaz/LNiTGtggu
XXE+G11tD6rm0BB9Nz1WtJqBRpMrfwnORaUNMZiaEdNgCVUbLW5k2cyYucTorFp39WXDHRB/Njpn
/YMbFIlBXBsA1CXIuAf29qqDT8wbBjitWlCtqXgPq+d1k/TVj9r8FE24OWDyxKvaLGOiv7AsQyPT
xyOpFdmGSKlypNUpZKSouCmPHHsfVN3XYl6jnmXGEPfcM8k5mGjrdaUfXTCGXkfYKDvY7r4MYBt9
9NcpsnF3le1dZNpBf2YG8jcQ75syz7GsFsHiJZen7NCojnZunYjgtgKsL6tEfJJ03RLBhls1UvPb
zmi3wVuPbHc4TNGkA0KmdgzVusdcTQ98ESIoGTVPSTekp+iaS8Gsfbnv6uATmlhLuc7yMsw9iP1f
kiEKOQ9DjosiRuJjSHxRlk8sQy0bvbJPu77psMGC6voNJJ9JB6P2BvGg9KXaqvh1xC2GdS1Owa+h
WycU8prPfFz8etOleEpvGuHUQOuUeuNAwiFtiOgwpNy5OmDZFU8oZrDFfbO9zhqh5CJsGER5oT1W
X/XcoQcqy2fu9qe5cdbBcfI5imrsL7NeDH+akbHyQQX6S5QRKPCFXMqMiwTUW07x7gFqwpyi3uBq
W7B6K8IEO8q2cRVM70xVV7vfvrv0whjxeAOdN2/llWKuf3o58hQ/VRHWP58qlyjPymfMVYUQb7uR
XF2Ey2d4U6nlBMK8OWd7cZoYA3EFVVVHdV70FvCnPnFgSU9hXsyg089Tu+Hd2a2NkeL/XHJh1EKB
G09qL6pBeF89Ooz2jz0g/WHfNHtUMv9ELY7TZoml7/Io6EfdMlyM0NK/CJ2CVBrj+HX3oW+fy2Fj
VxZ7gmxJ8PSl+aSMOeO8jJVOQAScAFKaetSMCjp/NGIDj/y/1+sQ51oWN54AMgLy08qiAz4GXECz
KGVVzVc2dXEefJuReDVfu1xTWYAUJSNIpAlcpTIxZBK3OZ2KbvA7cm4bgIc1sB5WtSY6jB7QNN3s
uOmdLMrUNkGPFI4oUfpt18872lW4XJLRTsgRUDkAuorP/lDbCYqnsfrD+jUXu6UJ18KU1rotC8Gy
0o5SnX3CIHIBeCDR6VOcVqPROpCiLRPAeEGboACn+lzZyUl4GXy47s1jITbmqivHe+2ilnEHdHoI
Bv6j4G74zHXMzrmIcK1fD8gVo9LFGzBYBbDPOCzXlhyF96hWCTnEfpf9CIPmnIBsQwCm9JfqTnsv
Q82ZwIa/6/QxILibYq5pG8AL+H0Q6NCL2EfrTTCyVhrfloj8KAqE+OapA9vPaG7mDjs0JOOwtPhk
EgEn4ykqC+CFli7ScvrYh1U6DFOqJe+rBxlMvEhAUuTzAQT2HpKiY+SCwIo6OeTY268zMU33FF6T
HEfOvJsIhinZW+iwRDj+E/yJodcUyLYt1WTPxnOYar5pS6tMInpbBeuBAiYwQ7CSRSpDFZLPpC2b
tTtdG5kDf6Sy3cvvtA/UrALJWoANd2EE8aYaUI0/rPCkvxsdvTCuvlxByBIuTSuMEpoiMTourmSf
uXteacbiVsy6hphwgH1DJ9ijyPuy9PgkYJEhV1avIWa8fJGX7q0/Yl86JzV5jrKzqmMf15YHRJ//
SpcBnBHuG68VjR0MVDohjQksh681m2ptMgwwgS4/wq1naHWfkNYxhAEiBKHiDm4R/1kUVbiTwjxN
jjThmgofWIVlDL3r978jGlmS+/lgnFAP3oZh6xFat53yvTGvg2jNAgoKnOBbnOOOPqQJMOPJXvIt
hE37WkHeyQJSmoMxWwkZmSU+ytCmxXZsd62nI6ma64jjA0vw9h0Fjmf4FAdO2UkL4vNDt+5bBcLK
lL400pJa9QjgVlWeFplfxfVszVazHr4/cvCgMZdoH4ShzgRENx2S5eYd9nF/BLek4YEfll+RuslV
yNIrO/q9R+AxfdIreqUc6tzYQNzF5Tfsqpybfk0qVgJ43sRUQgqD3ashEAmSSYGZq0GAINkrPd84
QmWAgseDmdYkibq+TWIJymeeRjDCvU3YDJpVLcHSxnnFW7u1DO1QkMboiFCv+uJB9mHZXN/3iCpy
Gk8olBQ3WfKKCyVpJfAQaoQd2YllHehU6UDelabwjweHrhS0MGoJculYgz1Vb2sVs6M9YhBl8dWV
4jkOu0ZKxntNjuCninSDedN1MQggKTNoIF5gzEVw8XOXEYkjAFzOwrc3VW+1UjwHPqlxRiaPiY3x
wfIZ/QmrTUaLhpTN/4cShb08fcNiNF3dfBfZOl0rgUKMnVFAUGVzr6AhEsYPm78VhcZdFvMnXbYk
jsltm8LY/FinN8PKPxngbavYgQ1FJ0zpE+RlDOLkV9gpSRNYBdQgt5NCcnbDZxVgph2kqaR1hkvb
q6RWR8gynluzSTFLTePxqvOr33Sa74iYkJb9Ozggx1njTwfc7f7+BT9x8tw3iOhz+C5eRYeNh+dt
QhkYfDD9PqSl6Ii8pLjCfwt1wJEkDJG850z5fRDph44Gt6JmyXcrA5EsouphceHEaIk+HDhwqskd
qrCHhVSEs8va28714pOOSPKKr2sS3XT7+OWIrQt219r3zA+JVKnDP31W++YgjmJLg1HPZSm4Cl/s
XKY72cPgN5epAaLBZujC+g1reo1Yai3QlEzBIJpVq3UyF9nBivN87QqeytCXRvLK/vmN152T4ySf
fjouKp65OzzLVovNX6YydhJh+cNjUCXPNNPsIqMNCqLGQY+uGH5yl8hkytj5uE0EnCrIGF8hhRXY
X8G9hfWhIv/v3R9tYwoT8RK9ToI5FWvctG6FJS0ciFXHb23/Sk8OIO23Mk/+LUj0E2BvEtBliald
TZ76XFZrvCV9KYTjmmPxjxEJnQcm5R2kxNYo0Pwhalf9YjaIF+XBgplsI0c04pWK3RXa3Jr44xHA
HZNDv0E9QNnr4rweZwupnReGp58mRnc/TqyAjsnb2ir7a5pLHyGUExdae9Sfd7gVoH8duBXUBQxy
lP2Ca8EaED1GsjsAVAVbn/PLkHa86uoKutHpsndlJM+qUPle9Vu2ZI/rrr3Od9CTpR773UqfCkvc
bnNToQUJvkwzp3sd4z8qjtiDwoXyYk0UeuvZM3EqGGl8O3LPcBJHjRGVNMZeUBQkUvchWWVCtyx+
oJb1K5tW4+H10MuXPFd4lZXirL61d5Wfd926HW1RZ7E3cfdzEk9rQIiDpt36qptkuYA7sUyZg83y
AI5VBy3xcu3ZvgcVbpQ5G6Mwf89rc2aBTlGXRJNESi6Ct7nFLX3U0ODXz5qq1/JAq9Cb77W7scgl
E5uXjnTdLmaXcPXQTEkur6fkehUtBmAqoKes3ztoalrZmntVyd8WFTieI6L6UFr9OEcsb8lAHAbh
h9lxqkemQ8K6QbQ5HC6ohXBXEXrvX0pN2hDvZIMLvhub4i4kxukqrVRhVZdsZQVi92Aiq1se/uJd
0QRYJ/VcmXSDvjfTuUzoyksdGdBtNj0P7IptwaG1CGzd6U2ZQmcciqm0t1zv9UNot74B9BFhA5PN
3NNjvOw6/q0lJD26G0G2nd5AobvBDNKAJr9mqbEYXcY9E7o0/tGwb9XhbNXDZk+Yd12+BNuAfn9z
kKIDN/OVq/q/UaVoT65/XC8lYPynlwNbPIfSzLYTyndXvHmNbOt9RtFSKeTEsEOKMxcXv/XBbcPA
LYhUeXRyOL2hq+FK3MSIbNOxQpaV0dSA7mb5XS6TNJbQFQjCX1EI36X1P0TqkNpbGBaBMe9fZUWT
1EFNtzsrCbCVsxj5RD/1ofzDLM1NT4+BfWg1hY5q+etkXa509QaftWwh3bUCk+/+nH91hD3m6Lvo
S/kDarMHwQHR/YhPQgkj4d2pR1d33+wL5GfUf5B2JEgRBUH+MHlC0JEhaWKKVkVDGv3EneVfVwa1
udJZ+Y0WHnAUeX4HpMaaxawkAp5YgmmWYmNfkFQH3PGlPjvN8Bk+rQzsyTwzYrZ9Hv+7NVc0J1zF
mrBAyPEcW25o4iBdyp+OU42jCgFlFWPh0JkM5Jqw4AK4VUt8NUttePOdkRTY4a0FfJplWZ1bsdhM
AsILmpiCtF/j5nKtNpoPURslEPtlYv1fFI70tGnvNdcgVFjIF9WsXnG4g9iQ3wZVzsopa//vKUQR
Nc5RrpjknCQRMCwc6mvNsDGCKBvlk6IMSHykrdtSnt3sKq8ZbFCXuRnIZoMi52AVpI4YytxZ3laQ
W5z9y4Ybxdfohhf8M09w57lk6V87CvxztI4Wl4nuVyHqFwDDKUlUS0+9IQ9d3d34qn8047Vse5zp
5O/cn7hkCJi9Vkq+kswvRjp/i8DiWfVbAFtyyU0e+huehKK8KNDvYEQOg/0D3+XX/2zkhHDn7Lis
ov149im8P92QQ8Mr17ZgUcIXrfWKhBYUYaDAYIZXtPr/xpae7qpQOgvZzd62HTng8QXFShuRn7Eg
NJA7kjuIcu3pskhAPQS6Bpo3HYKT5XtFyEwoXYxn2aVtUsDO7/PojdVF9fIEsHff4DSF2ON8NGBK
rUXugDNV3gjxwoaxio7sL7q2l9VhUGnWSpZyrOFt+qkv2qrJrwvt/4LwZUzxx7J+8C/mQV7ZIZqm
0wDd2DHuGi6YlM42KCxFGuRZ/4pqywWUjUfVTPS3v7HHAxa6XD5YJZtcyX8IWY9O+T5hOsh/1SyA
2FSp8/39PctwzH0g0Ew4pqmmCyfpCouv/7di/YQ76gIycaPSxresivTsh16ND+syvzOCw3ECZ9su
rEnoAcR6+XABXc5mi4OepNHXp5qyaiECDDGA0mGhE/NpAZI2Nkxlt7/+IigA8OBgp9rXVg1AD8RK
YoWBw27Y5J0muhN4vE/sGg9OqnC2ZSPk2mg7/f5luc3zAbld1OTSdcnEmd+ghClKyDsCiAVoz0pe
bh1os4VnR2mXvMLkxCnvq04zbJbYF3A6qdngmr9DknpRx9yn5dZC+xCJKoPCELFWWrCtFgHXXYzQ
JFLOI8PNYy3gjEdQTYmZ4PwEjpHODFUaz75YPXcBhYv5flYHmyDnQ+/h6PBmFKDBI1aluydDHcKu
+Uq+giHiBDDID45IGnjd+vjm6PBr4gvF6VZQwrYhar8oU6vUJlqcUxcDzTBJNxNgEvdNzTVlumjP
yAi9I6vmOWXvNaNdg+FjbNXxp8eON5xoXk6uVpw76YUB6DG98Y54hxtpAx2JnBH5/XK1ZUJR8q9z
jgozyJBpOJOUNCpbvjOxkRm4u1sLwbvwKLb8HTUjTJ4MQBl/QWzbdmfx/bTNFrdEAz6Z0n0fkHOT
HUnPDcqNKYxIFQCuw1mdSsSk4VqEi5abpEvVRBirOywH/56Y4zJ/qRk/yfeoDoxQYTbuXrh3nEmt
EYqx6kKlXfuFGMnG5ciFjbbmRRMYMGqsx5rDk4KAE+AORZbFTQ6ULaLB+6oLn5yMBXtYRDmoI7pr
FDvTYqeeJtPg9KvLKY3lXhDLcSfAeEgtYUfk3dl9SRQmLbcFhHx5h6YhkjRTIyEvVIQQ6NF1DXy4
g3rZzd9HqrBSdpjzitTJ0PB+Ip+toK6K5pt442KGNjDL9dRIDBxtsitQS4JZlajb1L9yn4hTTPdl
7UdSKGUWdJwGmfcoJHxKrxAEi1CuuHkNgLRsUSbC//dGr6FMnBd+wD+Ir4mZhCeGFFJ+X6ShQ472
8ciB6e3Hc+LVJJCStgFh50AoYHHIxYnF0nm2L6Ow35kAub/hqelLAW0aMd5Vvu8KQTmg4VLfspxa
V23Ap5+0AnNuzT0wB1QCaGLdTT22XXqVIAy9yIvW5weHUpKaDTSSdb0gqYN9GLM5WzkjgHD3Xn13
JAEis4cY84VrGFt1GHCqm0AxswqWzXkuqJxcb/u7hGLy4fIda+rtsM/HXBVtu8FUpelhMlFn+286
jmpaI4ItMEt4ATZwmBZBY9qEYCoTYfIEDxS7K/uWx53sfiw7hUJlYUMZvOHpELvqRw8ne2C9kxXr
ZDKsNjRpQYD3l60JZcvzcD9k6sqkgs/E7IfSGEiJp7l+GtndATEPXshP9XsUGq/xdrxE4EbZnNfY
MA3i1DtplBJUUlRS1Yi9RwklytVQ1ANImk6BR2XlNvKrbzx8AzDda5qszA4hwDRYt1/mmoRAdz8i
fQRXcAZ5Gukhf2kJsaFJZ9oz0mmK/XwMQfw2zKPS/1KfDMw0hEjqv+C6r/Xs0zI/R2c4uZXXSutt
qlRcQmFn2W0Nbp5fGsmrPL5QYhL6OJpH9T4AwkFp203k8qMriuOnGkMBr57+fbVNk9d/w2SgOhTx
/jN6Mzt+uOtKvu8LtCHavB/8FdwzS4ZMxp+EvmydpJcdLFIAmqwfaGphBeiVngWxNZ5mJGC7C2f1
OSkI1uz5VzLLpVdTK3l9yLN3IcTI0CMPxoaXn/oyxcsJzTDtrnD7XsmCar3aXzJe2s2dSNKUcHq5
bo2yBHVgmAMvny8HXn8hHjZPbydZBFheAWcJw80uuLap5Upl4QSDfuHnjjORhjEx0g/scNqPXksP
WA5nWoAHCZYkJiYvZNFK1KNmVXnD2fALAghNfd3nS1h1WCbwhE0+Xz74b3GU+aYyT3nziXVOP21a
mJQzTuv02AI0cablXa9x6VMnA1xUGvlDU09oW4hJsjVsoObXGTodEEZAlNb8EIpYOPp0LTYVyX3C
V6lMCr2tnc+8iO/z0eBapk6k3iBLf1bxztlh8MaKAy6eLn1+ZS5Qrm4v3J4KZlnjGe2Q8M10KE6I
c+b1NUm4XyEpJTu+oBAeMw43ICMm2CeW33F3HBLycBtwFOpC+2BV6fdwQOmGVEnEUqKL7O5KsbEs
pbZIpNZ1F8ebqwLd3j1gbLsoIrTTzTEKddncfRxRrB+2dd9lhAonh8NFm0EDm6VYS9arx36GEK5J
fNJo9fNHsz2xFZ6sV5hfEeCBFcRZAsQUI9+746jOS6qv245+Qh/KWzzmWZYnLtnwVQTozRl08kLD
ErSoPkfpXup/Z5To3E3qn3gv7hjB+vsf1tINIa1WdcJk0jjm6M0l0m6fF7eOFmOjq0QyWdsfNgEd
YNMZ1jvJhMP4mCZuiKBpmlHzRoBYJC0MrWXViNpB2BVXwlR87qwjhqOmc5rJqdVFNuoMNR9D5D27
FHbvwK5py8bPHsspZ2Pac/oh/zDSi/+M3BkowO0JegatiD/XsA2Caa8e8sMMWE94r17iugKnstzh
Oqvh2tc9zZuhDkAlVXd/AdgcrcYIr7lo7glO1VlMao57dQTW4QroGM9V/3eAdfubzoE8avstyXdv
SAQjb4B+jVtjBJzh1zwNnctI53s0qRwm80HTOASrJnNtA4eouJU1QHbIe2zISIlxl3GpSWPTFPXC
4c+6fa2/QNA8th3KTOtSDPH6OpWYsS2PyPf5tZCudQuB3t8z7GddphZNala6C0/cDLGf26LHLf44
rIPrM8bizPB57hy/unEoS9aE4HJq4DSVTDG8aTwRmtWPY5nynff58pwthtr+vMmgxKRSKmBXDt0C
xuY0qiWteEdhb8eH+CjIy6MK4eSI3klhHugfk3SjDbi1U1UTRGon90uFT183ng/9CiicW3Q5hchK
gpYX+RF4cCnjT08AgBO59I3ppnUWfK8B8JvfKBkFx8pZuwrzIFYY05yXWeRGv1oUk5GJ15hfyRZX
eXZxwGyjtYps2hjpGNSz/MtC6RRvT5PnJuT/UycU43vasXelprkwmOERccIOhdpTPo+q/B/IoIOu
9PHjRh27cVBvxdORLnacm7KDV4TVgyxtpj1XnwwmxBdFp1Q5w+iBiLqNAuQ0b22jaEPHMurrus0U
rPjXTySxHLRhoyP4iaPLp0Pg8JW58fnzrHgS1b2mXF2UWXhn2VS0H6OO0hJ8S04b/C8tZlREvQ9+
OimCiJULR5pOwYGKtvreefaFk3J8tF5p0jkEaLSwRGQRAjcD1dTMDLSRC1xGvQeTUqLcuDslB8VZ
vsqYl/FG1L9CpcR9YWPBRMLazf+v+QV76tRSiNGhqBj6VypXWB0AGJX2rnyhzyy2ZTcvqR9ok7wT
YZPZs1ictMefLPMcxJbk8V7xwmYwiKXGPf9Zr8HBRO0Vi4lgd1u0k9rgBjxsXdCpcacizWZ4YFOc
7ImdcbPolx9atxJ7egZuXJcjLyicN030oFpTXtry23JIrcHkE6FnMh6fbNhgfk5VLVpelsKZiqaR
tDOehyHtkbYr0MQZ2kITiLN7Jj+OioyggBZZiMtPQ/CVksDCRySWCCvHfUnPOBIvodetqALYVdYO
r4lgNvIMEfm8weE5mDuqsxJlsg1u9Ji9bHQ1atKitYSI1uIqfZ58/J+iVvx2UMqKmSkKOGw2J+vP
rts4RLlbr7ViPZgqG+v2TjDAk/GARbV3KPCqKTaDA/DnrRMbP1svup+zzQG/x3IXnfchW1Xp8TYl
rX1YgZrwAoOo8x2nR7gP2rvggWbWoPgbeYwOQl78rh5pUIPHQM8aMzifGSz/deFQP+ZWuevxFQ5+
Ed9DNxHeg4JrIKfJprh7Up9KJV9et5t2Pm1fpF0EcG526IkwDUJdHyrtx2GP/v1CsDrDIdcduzei
adJ1MIQ64GuliJtmYNf+iy2hrMqPcJQXB84VMFK2RGVax55GEKSi7CLvHTt/VVjDTK1UJkn12Bcd
2LWG3VY2uw3Qd7Ilp8c3x3ztNw+K2xNQtjwDSlZp1shfaXt9Hq1VejlUWtjApdgRAomvo66kUort
hFmC505c9xepn3cBC75/mghDk/Oxp9oIdM5bHlHMfLT2LgBrnHSRlnao6mxGC/sn9ldDPywx19rd
BiFNZcEhuiWiDdyV4qVZNLPP3rC0ByArNPI7WMIX5F7wx74e3pks6eQfP7St6KMgaL/G5zFXVMiu
5vBOI/kcrbYiWV5d+n5EPrYGH88fWPzD8u1uQDZwtlItOwqNSP+91DK5LjgjEhQH+yD3nzpAkWO4
OKicJ/b7Wn87h6sBBdZ2M+nNvQ12zOD8Ebuwg7Rs52bnQCznW9PvsYqBumjPyt0367QKDrhVMcfF
MOrAJqO2/jwKchHQFD9U5ezWX7jYMjmuwJ466tvoVEtHphAMzcwb6RYVm6UUczl77xa2cia923+I
a4DyI62BGCYNFctv92XlpuPYMZ+bOQqGB8qYbTha1z2mv0HLDchoqLrfG4Uby1oX17gbm3CMRt/p
PdoGKZD/80cfA/fp6QmfaP3nmfboI6iajzRRZv3wrv63vXe6bAuTtgrboFMN0nKYWelUdg2+0gcp
JkirJlDhgXxahRFdcGQreVDsDJbaJJItdJI+yhkyg5aYWJ2rE6XiGbUaUBp7LcTcNt52KNrfQ94J
FbrVc7eC4JTM/wg2AG8DMe+yiiaNWBAXlbYQ7wLav+Ocew3jdveJxyVI8paUhvYoePP16eP4qtRN
KEHs1lxpyac4EgQMV3ABuq/rlHCIwW2jtWuMRtUF84iX+xijru8y2jYdHyUq2wl/hCinsHKe3B97
TZI1ev4/uspOdazWEQ66aZoIdoxy05PZsTel2shaEogSMjFzKaBlF7C74yIBHu4G/0ZzRJ7QMWWm
T8RM4E6Y8C/NHqRB1j6qhLlCwipjyVoNRN+wFJGngmeMX+SSmiXxcu0zpFSQfs8LYElrL40zAVFv
Z/c33VTmFAAET66K4FnXoa0szrhPDKI1Nd5ko5FX8+qT8/wXrvUSomnVT/A0S8tZrMUuwGXeRhmo
phiI2tGw9l2lZ7c+pwSUCW+47K3oe8bUCIMjLCK9QdlTDe0/E3rTIrTwLKTsUt5ZoDeZreHMqQPa
kXix+GST2KPPo6xD43YSfhd+awSLJzGpyS9/+PUVyQUrqdnsVfeFxqZAwjJgxfs/uzhY6hZHa9Ez
TU7BfGwG1/r04vAzFaa3BLPrQgavjj2SSqbay1woVIlYq2OGCTAAXbNXcE0U0JOlz+xMxhcFXzZ4
ZB+FsxEGCjifW0PiBBvUD1mRd/+7YxGzuqmngHyxE96FM3aMvcoGIXsEusXYJEA0vW6KRgXo0mcY
PNUfRE4CRtphBSepnQrfyix2MGQ/ah5CD7kCK1WH0PrCdWvp930Um2mJR+TxXtd1nWgM97YLzQP3
YY3JkCj/ydLOpkhYZZOkcCXjbvgPKOskMsyaUh6XiHxKGLT37/6d6vokRz4zuwe5Q2I7lERQbNNO
axqtmjf/2TCUUj6KIL4n5HXJEfcG86MzHtc212AGHW3NasMEPo+c5bVET7Bj9mNlHDlhV5RanQ3t
PM9ksleZSWhzCQsUA835631n7oggu9ik2H4EEidyZ4PzsK4LHIlfOdZCMe6h4GRwS6nqnRudsg5U
zL/9tw6CuGgDpsUo9W7vmEz+Wga5rntjsj6VSw+RQdpAmjL7cDtzC7HaaBPR5F147r3qyYhca1Sr
8NQ6FTLE7ZrSHBj+Z0LTrhQMF/BxWQ5I8hovGsRC9gvEPk6f93S6q0v4rT+Yx7hD2MIL1nVHE9mr
Ak4hPCb3i1h0kj/vVRYYHVtaeitlvjm7XJD2x6MG6JRYociD8+vAA87nZG70r7Ed1FRa9qOjaiUI
vP1V9cjTvwj+Jy0O/XYYtmEANfojPYhQtu65MsbeqKfp4J0T5M89ibiXFC+Qvqxr1ZE40HNDvroz
ZJSRWUKO3ZqPLb4pPHCpU64/nrjph/iCfqHmzP3LBQ1JHoYoCxM8xsX4GLapfSFR5w/+v4L6ueAO
s0YtZZfss7bfHet5N+/zBdt6bODAnELLPSrEvEJ9gLBg1xxdD8cp4AKC64GNdOqgZVXRp6WZQdnq
jxYWeVwikftStcGUpqVE4X6vukvXLwVvasAeLFMQDKUL2cLXL9XcubBff37PTrq7JA6+UYAoLj4D
xLCoyUuZCV++CHXlFUeo6sJRrPoowfi6xUAqms5Jx3vQ7ch1QWMnPJ3owktHXDQOPEHWdzTAknF1
CExDtMlPWQc26HQimCW94/eaop9BNLA76JqTBYTBxkonCztF0wpsKx4CJlQQnRthQsRwbyL3QkX0
mDSmQB43RiTWq76MGTQVHy1hPZxyVRJ0UwqONcIHPesl/eSPhZh0lCTDLX+pUMjna59Xg/jDuLjT
tE+0uDHAN6t4w5Z9YxzOqT3wI45F1N5nJRmWMIp1nzpEC25XF3qx9P65lbqwzHB42//o7E4GerTy
mfYf5nmLkCqpbh43yP2zxPGdg1UvqoEooRL8+SZIBM20CshzMDEVuyu1tfekN99mHSe/qTSH1z11
Vm12CHksgdoH6FN4q79fC9CRIirAzX0bJMjAbTOwfiOz+XaA4KUZ5J/2MX3Up64VvcGlJVfAx+bV
OcLSyMSWxiN01/g74hKAWB5iWhIoM8ccq+vXvPWJXm9np8K8j4vXHIHEX/pRmEyDcrEfKC2nqb6G
qUqvtyfgLGMRo4dhMu6yJXhvxZPyECxK3m+SmdDoYRXwMFgyYMbFuQg7/RK4NzmraiLpI+LnC/IR
p9OAjWZuQNiffwCCDpm+0lmikGo8/VOjXVyjq9cqPqH9klc7T5OFjc9uytYyNs6Im8PU7xutUXYk
RUyhFqP8CsLMiF3DFhdsaUv6LcBBSjXZgGQKLJwPNsEFX2ZYnI54vw4QgaCFkTNpEAGM9cazEDe5
qPOYr7I63ts9jwxHt33O6/Qun0aHzWb6rs2aOqkV8NNcblVXvxJd5cP2/G5ReJn6WkvFf6Mhw8uq
YCQgQWeyki7litGaVUQ37kclRaBIVm1gEq+v8xdeWwdL/2tME91NcWyq95qRfUwFG1XHojml9r8q
W4qSnd/JCLN8/ekgyOiv6xdTKWAhVdvKLIJ/37veWJmqVbFOKIsO8cqM1321FqoyGKMfjEAsGZkX
ug5pH4D//lRKghznDOUD5WSu8FS6bpUVIGzObN9lVv+AIJLofXVQqdajL1dvJeUkDbY1rdHE6i8f
MJj1zoha3sk9VJZl/R1k3zppcHOwWovaaKXStyLSmaiWsHXB5F4zRCi6dGgh5KQzQxIGgAHkVJiB
AoNf0i7Qjk5axkgFsTcg8k2FRy1KeCz7apVMgJgbDSWCKgZMW/fgPVGzZhl9BCYWRC9Aw1aOGuaH
gFGHMjgZrYaojjqaeCoavy8nbP49DceiPwiVk4Yd5v1TlHMG9rPXOO0l2M63H2TpuiSJWJS986Q0
KfPVFqUq/kYCiCUaAzQuBXnffxerYfe0Zg3auzMStszQ1AuxZ0qXDlToEBsjA189ZooLo1Cdg/65
6X407hxeuA6aPHlFn4IwrrPUr6OVFWyVqMszMl67vrtrKkqVTkn7rJEuiTiS9K53udt7IJBtAWkM
zrKs05x7OIhb2P07I6iwf4cUjl62AFKSuzA9LrxN4N2sQhl7LPOSjRJQvqn8BTg6n76KTWN29XX0
e50I26+exAM3Ag8kDYczWV3Vz07dkCn+4aAOzHqQ3VPu0g5kHv6a/FMUXN2o/kVckkeFqjxzynNU
IAnnE3DXGns++/syLDaEUVY+1KBuc61+nE0d6VBtjkD4bhYvP+KlJXzMh360RXo1O/SoB7go3SU9
H4IATVDLu739JQc5eoLnonUGCZh2rCDphTjxziZL7UCGK7iSzE8971gqWDZjUU8gPfNYEsimRk3s
um5gjxR8iegXomRAIigrZFu4tpWl51JOa9WhQ6O2LMV3IrK22OAGAIZzxoZm8nHQ9xexh3HcpVTi
PUwD/8iAoAhrSMemNHtZa0MjEbES8BeXkEBFEmQneKCWrfZ9rwjY7XNl5b/hnuGpej72ZQcnPzpE
B1XSe+WZSjrpdarD8ckwz33BWlxLFx/kL//0rxJxte7k9Yq1XeSWzfuODvxpSp5a23CZa2stkkib
XIV9vrqOxrB7GrTHiOnpvl9axgyHikhxNAQANyN+EIByjyIGMwrVag+pjoqavP9V6drGDCzyzwZM
3EB7kJnjvVdY+pl3LatsOou7g3yDZrSVzV4dJBQFI5cMoTogylaCCrkxe/+es0+tNP5IrXMRGlLD
NqD+c11PvAt6nKZ1BhZd4hxxdXH3MOY1aQhdzj3OSd18GHfBpyrMjMg+12amrH/dYE2AhL2Cwt9L
Qy0p5uUWwhq8958x0EK2RKVVW1OQwrQxUxI7Hvw9tdMpQ3IAkfDtdq4knrPvMsP93LSKAQLmpR/r
F0S1sthm+CglrccqM4eU5mwOYczGa2jUAO++77HsXM4xwsGRc6v4BNt7uZr06/jYszKQVeen2mXb
N4oJUJfwiRlE9TXfHQyI4F0Abi/mxI+POPWMCbv+0xEDpLgR2ikar6nrigqBWmppGdunXuz/XkjW
S4vsZbaGfGv7La9Co5EtvqEr0MBiwtCt6CNmfJldGjsC1N5O017HqTF/CQnJW5THmdvhk79tOkS6
klsgZoa3MeHHiDh/rJtS5/JxrQCeuII6eGuXswHghy3K4m8jPsNF8T2myC1gv3n98OZsFXVl46vI
IgDtjNccxpqMCYm9IW1RbzF3k0RkqwJvHC0SFwPMM1p4cxNwFIWMyeAae+EnMeXl+gsjgABdS0Um
nDCT97PhTx6iZ2BdoUFJBHc4DXmnPxHx6Be97QEy24iK9uzJ5/gQXjhmM+zpDXgNWd6f3bYQJTw/
OxHkibRaS0AoT2ZIyLrxNEj4zpeepabXvooxsX4ga3YclBRikMITonPyESj9XjKmzIqXrLPezrqh
pR3GI7/HxIzl7mOaZZNi4if/wKW8+nZfz9idhXZcFEyOFgHiMuYGBCL+s4c18abOz6XyvR20Y4KH
DGecBjCgAr8j70TNTR4e06zkIxVAtLHcFo7dWxSUrvntEgQFg6WrS8PphRK0fYr9LmJyGFx1SDmF
o2/IQAEnX7G4yMrv8879Kbr+q18Dh44nB7RIu8K6ZvagPs13ZHWSol1l0OKmnwnLlNyErqgdzCJG
PM3RDikBcLnouWcQyZKeyopqiRF8e78/tOeolAmPpd7NI44F90Ke3P5CVCmtUEMzW0o02s1azNqo
nuDk60nUwO1CYMEf+NV6U67dve2BKxcYCzr2+bv2KbeKvZeMleg9DxIeT+hKEPbF7tUbRDTqTyjq
Eo6bH74zQEGvk0Af5p8JDANpY9LJIb5wrYlE+R8QxJ0vvM6LdBMQ4/38jbjFjoYfAqtSJIJ5yYdZ
hkSIrtCNpvjVYalyYW5tomZJeMeIce1mo0jyUXIoYPohzxzqSb6yVSxJXgYONGrAfK/DbvKEEC5Z
3rH6fElkODGNMcCNQQQPelCNHC4HTB7P+GXqZBljSm8yTSWJyumS0BeUWBUwf/pk1Qve77x5Vil2
XooyVKcdpwKV8UZLSvsUBjXJDqq5LYlPESf3Qx7J01V55BxDvGNKr6LN3vEM7tse42cRvKpdM50h
9NsSDdNfZgIoRjzL/R7i7ZwAQtzJ3AI1/BLCs78P5TKmMYVy3iboahQHb6ChlryHpVZC1nsyvqdP
XE+moSC9fb10xApfoh+4ZzEOqiRWCYXwm3ISGj0eH4K1txzOGB9asTuJulSyagT0O1LTTFCrigW3
cy5kM9QEtNPVBnw91/Elkm+IoVcM86SXMiIbXwyaLYxl5d+643a/E+u1rIIhoAE6xi5GwN8xFDWG
BSJIwzfVroIjibxYbEXULjSXED1mfWHHfc29wsqx4W0YmgcjUYqg9VPPncOU14agIGuWMtjCCNfa
OTNJ3qKmRqz+dEV72tob0mI+6sow3RWXmYUbp/jffGwwFx/UV9z2qT49Xouie758gArFMGVlZECv
U7aquT33H8EcCszDII3st0hO6DW7rY8aK+ln0765TsvDK+JKhF6dGmwA32SBbUpe3oB/nvAEHuYx
XfcbzH3ZDVQPbt61q/33A20dLLkWgCm7SLW7Uc9BkFkZ2Ah3q4c1p0XQc4DBAbMFjH89ZKbEHPrh
zgNQWrE++nWcPA1T5i/O0N9OMY0iRAVYLJAYFHqIRu2IHDEA+V8AT8PUdFeQ53xBn/6sKg80LJ5V
3zoAdiJBkwQmlaiO/ai9sPUNTJr1+ZD4bzSXxs8MB8dN7kcGjHN7PQcvypfW41V5+e+zYJMnORZL
Xg7fMvi4Qh/2I9VdTXGXYOqClhaB088/K48xW5DugXIqy+oFePTvqjRz8lzqJ8W8cryvecHe7EGP
GeczYNc6sn1PP5YOe3FsteF3PmEmN+i1vR9qux3UDPBzO4Ek7/Yo9OkT/nrpfDBQdDqv4XLLKfw2
/q2mhnbI7BpYssWX0Xk4eFttikdwxr5T9aHuA6QZ1h/jU5m+xImhMVWQRTCi+/2YzVYIbsm0DYgR
ulS08EQPu5qIuRSy/UcOsQlKoG0IuDHX36QQ965QG/dk2VPiICdDrfneQ2f9Hfclq7ycenOiMFU3
FMYOec1OSfkwdaFWthABC9ybahjT/czgx93iRTu0/W53n98Yq6k0B4pud9m7ZCbYlJN40iGmNZjr
ptxafnGAMMIwHpdMR6UUkw92kyPdLORgZKWOWGypIwp+lNEa1P7d1N/L2/t6orv0YevqmyruZEDO
0TzJ2pYUegO1MmaxX3pwihFR+0FM4mxvKHeDsAEIPjSlGiLU2tclKiXwpKFSmPEyaQ9j/zFUXZVb
We5RBBZoRDhC58oTEJMSSCuZxOuC6whPw2IlYlPbBBxlQ62hmbsd/kDn+sob4nMk6V1bDk1sKR/+
/D//GtyZ0Uxzxw9VI2fQx+nqzG1T1XHcxx1Md+o4aX1W9f46x4/b5gtsI3CPUPGRyt0Rmn616KnC
DFAWVAdJdDHV52ZgUXZd2e/cx6osB7tmWPaTU4LwVN/lLMIv3jjpekYdjf8kZPwGaNYwaz/3CSR/
+P6FQOyftlYSOGPjEWdVmwBspChzi77ldlSG+I5stdqpVnJjiTW/nwJxA/o0gwGgqGJLOUHbHzG+
4GYpNNZsHGiii9Wy6gW6VotfvtQeLeV/UJXIouTefjYz10rNZHltux7/AtcYH4v4rQdFMMCzKewe
sX1APIz+If4REnq12OcQIA76JxpIu4O3Y55nhzvX/LAeaNUNu0Gp3jPgR7mYkDdtPLyhvpF00foL
kpW2RFjDMownOlLVbD4OJYR9mL/AhUc4L+JrkMqYjJbopN/m8m7uA0XGT6Inz+j9ptYSAQL2jOUz
hz2rLVqErTR+T8My6OouehU5n5XO0GZ3HSyivsqEeKsjpJRGm+Kcsx9YBbkL4bs2xzObT9c0WrOY
a/04haDg9JMRuydFwu02xzneYOLWnkICtP5WCVtj2b2ar/tpsFUC/4MFow/lxTQM3rBIlWS/zLU3
7vnrxmADed/Nw5B2RqUNJ1E1Fs7q9ppO5M23M/j50JMtTFShxAhylrDpHhiPaPCOl/Q5hH+1PgfH
M3sq5pBI8ye9kTjU8t5pgIuzsUmjnIo6JWj1/UV/D0OVUulvqs6kT0qijsBvnAfVoEewgjuEUpVy
RhpArcjd4Mwn6mkPWpzA1cWxPw7Zr/nsLck4yPdSPSYyT+V/Kkj6WLbg42IjZrVe5i8UyQBV7nwB
xgG7B3LMsONmQO4TCieAKNxjUKYn/K2Wv7c/Nigguor2A9FsasXTSw8tEYAFqQIwSgZFPKNNIGfu
RyVinlaCVUfhFXsEfJafxfM4DH8EB+COEBaPJBH0Zu7tZNr4UI5s3I2tS0J94p8RnMpt7kbuB2lp
MSDgihznhb9GxgI7Gfq2ZIJW+FfLzGlUrt2D+N+kduikm5zUyY9eNJ7JD54a5QL71xt1H+ZaCCa+
OwiVM+jOqjqjYdjrFgSRMo35CctdD30USnZDCpIJY95ppDQCk45Pv3dHSPbPlQR6B3oYr+jiETNp
HTbgPc7wRRIpk4QxFtmW4lKIiKrL6gHOCzz0BGdCtzn1XcJ9HRsQjp7CFmA35LVL1D6yJ4H/a1k1
wdFjdjW/6K/GpP4GdqIEUQBjtPxXFrdWhUmbvX7RB7yg1tfvrayPK5DyiEMIPgOGysscMQ7+kejJ
o0M8WpspcjrjLMWZ+uVneZA/pCLgCf7EikEd3TdLUrui/ojpY+Um99dQ7eMQzILbxM+hUa1h/Qv4
7jH+YKfUaNEcFwdIPNBF7yrBOBGydld/cLKW1n9nXZSipyzREHglFBLfq8TL3uwxr5k2X928FMiJ
AiPtwmUAAm9slH1Rg4yP+hG0FYgoCR3hcsUUt9fLZRs3NGJJ7E/+r28vTIbKIvwke2mMc6OCjVDh
q9OgX1o4bbXBf/FiUCliADSZ32psJFBHG/0HSyhJi1BkG8rfjW/OEhmO+4VvQmAFnkTj7XK89FEB
0GPE5QVk7ptWL1HLOcbC74ukJbljuPYks/v3WG9Lh01Yq4eIjD08jpnFm3LABJWZu5Rh2nAiS/aR
CMGkO1EUx9mOnYodUHGXwCgqlAn6fiAwpJZZ+XynU91gGler3qz8/A72gkEJ5J7UWgBJ6S1U07xK
8fhJk8zr46KXAfggpTCRkOuz/YDpr5fHKEMcJ+6iDTrlJCuOZffKov7avuPmUyZHL2+4pyLITWFZ
TnfOMZYih+3VrwQHNf6ijHobsW10/CvjN3lDmOGjcuvZ+pUOd4P7uJ1tckGWUbWRVnAdOoKDWxku
Y3KbzIe2CO0WHiEIXxj/YZSrtbh3iLhQvBc11y0g/X+IwSrjXRCx7lKILMwgfID0b96yGLLGhYWI
80wZZvCBOH1+PU+LxkFC5mtxBbSQHUY0szzCXP7sfS8LBkj6dT5p6RabaXJ22UtCV1beGnyw+Q6h
Kr/hU49GHKQvFlsRxIOYmtVFNfNaLDXzavLifB5TqnBceJNG7+/hU2ux81tbKvP/0tAr1lwvOM+8
sPEeS2wBZnEGjEaDzOonKMEdkXwqKFVC1YxY4EYAJWZgBKWxzCZVeRZ2ruPDQzXz6x8t38tikqTk
y5GEgNkOJK66fZp8M6BA2pKRK/fE+6bs/gLxmOzu0UTgJYIfbZfV2eDyhtCCvK6e+VyigDeg2dQV
17MCx9KoThM1OCv2yNbDRZjOrWte3mp3krlFCaC1/6s9mJVIros4NP/V82IgpniwffFIiiGrqFJN
FUTs1Yuul2l7auGdf/jcNhhvbTrZHN8C6jvMLowzR5IOvm1KXWhI7ViPbZNFlwyUjijd+5YOaBKr
QmKx8//nyKVJ4+eFpQKmAdP6VDDW2JnehFQ2htZp+s9NDZ+XX84ZM0FcKyu6DQf1Lr3L+y/CKfsS
5AUTKfForxKuH2H77XcE9HTbFEbCIPjfBiQwLawqTUUbmeU/B01adk7OyuxNwDeZF2cd09ihyOcS
ED5c3jByXjBGnpnVmQdl4Jw+5f6ZSeUK5LNTgFNOub4aZt8UFieaawbQDsQvVYnyJiGcWSP+20a9
jcA6DW44aZKXc+63ukdBF+OvO7386JkKI7E1Lo4ob0oVu0FhVmKZzZKd8LEqkY/Njv3ngG8r8L2x
uSRf/tbDF1MXs7rnlKWVDxpQDiAmYuNlGcwkJkyDRZuR7uJ/dBrF22EQI7ROiIJE63pt/b1L4Sf8
KVUtqQdROhlsqDJXc6TV0sjuBFN2JMfRuI8Olud6dOn68jrN/DC9ad31CUahPwXxMiQ2fHOANEnG
iNGZ6eKEYR/UETd+Yqj2BdnA3tyIraZG5/9cC7UfuiqJlhQhY0oRjDEs764ysruDxyXcqIVsYNOL
5dznltqpP+JE7uKKujTAeyFgORXQI8U5pNksqscqlufzEk60ORSfBM983L3cokIfCpGEsTK5NgOD
COkI7xQhQgfhnPnBefQbydm6qcZwkZ7diukevhy/WnRBNRw9SeCWr/cERrBag0uGO4KEXJJlq16l
JSTEbGqxGYINItezIXB3+NZ0Q52H1jJj1xHeyMJxOxMR0DJ5mS9JnWDrlC4ZSsPfjy/8Ve4IkIl8
MmjsJ5w7wzl6rw+eItcDjJdXBUx8DiHu7CZ/nZ+FWMjtZAhn2NV7cDcQl0xO18UHdphITfK9pK1V
ipRYMZ4PJ/gs6vx6asECDblAl9xY69nKJmqeAz3T21XZUbuKfp3kuMRZ0MyVvAIV6L9vcq/8qa4d
aw2uVQBw/XStwdIUCIK5KE87Eb3olnkiHrqrYnrkCjo7ggk8jDiwq08iWaA1GsFGf5fCDJYN3w8R
V6vyfv+KbqPvz1km792q/Qm6/9xdF7HMAZ4TJeH8JSGEZJ4ZSzbrjZBZRrEsOmYfpd1lbub+F2v/
PqvKluwgCO5MBZ8eKpGsoAaBIckX/nsL48crJbzNuHyw783Z4HG4sWdsQg28EHG8Du0+yWTRn0Hg
V2MKRwOfhddYs7Yh36U/9I/xwRhqsUtRj/f5lVjDfVQODfJJazOXAn7osc3/QovVjDf1HYpId6Jp
JsXZeaupJRVjCgTLB3sbd/9Q+e8d+Ujho3/65EbkacCkLANxFhOuwTYeij3OaDBfDV6rmUoq0IXm
gnY7Q8pwJjJL3r4IiO8vS6lQCi3/RXrnt+7Bif6PBq2cDDjhZT9TWC++SqF5M0PDwdO8DI822Sf1
RctD8DOfrQotGYrSsfQGb0GbLFomeyym7S1JhktAOMCekpFcUfcg8emTk/ohJZo7BJm0M2y8gD85
oFtGhd8bjg1hnMJgWeFiGtv+cy/XX4sHjlIFwrPJIBgIkSpeKT6I2IyLKcdraADUnIvyq4sTFg3N
eNlTJ5+FRz4OwcvSNgQtv97URmXA/ejVJuPOwchatfCk1e1Zfb7YFho0Fbtg+4uLwuAc8rwTXCiO
Fsh/tVFSP808GslSorzWV5oSVjAl+bbkmdn3nLZ49GT+MMdd15CjTIX5MBztP4Zxk7gzHZuxBZLg
ZC+TyXFC+/kZbhQTUl37GXU7U14DmAOA1nvm9CWfJy1hPJNodBTnX0kJrklQ+TZUz9NYLAmW81mB
tI5Y6KSVnBYn+XQT/fpfheAvzfQ7WQNre6ieMEKMrfkWTtgeop3bACDiUOLCgQCtgb+z5Q63miH+
T8OshurR2mOkRTOc6+fga6NP1E5GZCUJ7DS1hFB6MCdCBxaVOIuiEPRR2hvEsovbFQjG/P39KvYk
Q60poqCQUuJWhL2oGdukf1oq+Eu98R1eXkXcHEcyA20l0ZnYE7dX7L1OMOF9J8Y63ZtPxdVeEYxP
grW74Qf/589AVCzbQnCwIgGBVLyysKWCjYYvmwxhYZnil2HR9HMcRPr5wgyu+K/OEX9hKQQxfFvt
B9n53skKJQEQHCIMXYddRbJpwO88RXyNxEO0UXSNct1ytBRtqad8zSl4af/tdJLSprYouqlvq14e
t6YYXtFGAsuJkucMhDySwEzmsrCXnyoXzsgX+PyBWdC15OX50TqNQX1K170D2xlqtpRUvXDUxYwF
vkppxwSvQwaQiIqf2FniUdLvrhxS1TO4d/jVTXb2Y6kCkCJuUX8AZH9UjzjwXNKpsK6smEHEx1JH
jwklLfnYWZDpzliTqghbxluO4DDYYP81YiyPuvFPyGE7aFpuInx4J3dYMQMBJBPEpO9n6Nh79SC/
HiU/U4ic0rkAy4OKYMmDY2luC6jamXi1XtdqH9cGED7cXvhOK5SNaaSWS+TzarHVpZ6nqMutqj+a
tYiwayNkPGZw1UgyzYRTcfdZc1R2vbviYpQdGwaz+ueD9NeJ5gsRdquAG7XNmKstZP9vb0/29aBw
BvkwSXnKVR+yGMDPloyg4cve8+R4+s/jM3ediBYbSIewQAQ5pJ1FLDy7pI7jTPIAFOrQMRUAMh8R
9QC1ML5rcpfVva6kwyWHSN5/TMGcF867dK0A5hAcfMRILrtWJT+R8KU3xXZETR6KHzsyHKTxXrXs
MDETG6TM7IXqDbpmeIz/SSI0JDviwWvumzufuyB3etTVuPBupLZAcBeE9RSTIOPT5esFBkgb9CRr
pVDjT4SD2IWOgNF1RSUAwnQZaP7PYun+f8kKpCunmm71CUInVwvWTQ/3XAdiYVAusHcIJ3iuzfp+
z+9O00KypyXimacPrMIouKkApzvpl9S8apFStz0yey5GaaGp4G0zOHqWz2kHTetO6KKk/lVG2Yxr
7x1hdt2QxCaiX13yRlFAZwM574aLHr+cLVHoAU6Eh1pE4kJP06EqzxZzWkyBnBbMQ466hMmFrA4u
kHHOM0z1HQQRhnb9YyjtppkTM7qAki5skaJWS481A70bSuDTAOpJFv6Ff0UFFxMRFJHHwpztiGhh
imtiXf5rppiX6FLNrEnbJwtq8Q8MerwwuIioElMczUtp8naM6gh8HMzOe9HcFB34Rp63Rva9SAjl
wn1SYf2umV4gZPv1y9Y673hNHxiyjzVqYElICGlJzGMGSMIusruYJRlOFHj9L2fUnhx0EZj6sSc/
6PvAppeOTsjVyJItzJAE8y5kIpEaxTGiWVAcdF6OlF1Op2aJKRx1xeHl5E0lKnicPQFgx+6y0EYq
Bf1v7FTwEeXikAt/wKxq/9P9tKV+cZex7kj/I93fPB5DecJi/C0YWa2NHaGDxNjoFe5ZMOfjhprM
/Py4uSVNSFNv3hWIWhz4nKeTAeTEzZR1MstEvv6fkTsYYV5bOk805AVvDd0q/k9F4giawDNyjwzH
yShRkV5GWfmYdkJb0dk0QwoS5gFY5aLrK6JYLMmrXY7fd94LO6rdYS27W1HSS57bwJ3WrZxac3f5
ec45uoaVAmrf1Q4twGJfok18RqYX4BdJZ8i5T8VHYn/8nrZxaogEqjR3LVeqnMdJB3y6CXlP9o8J
LRPrN79w19+zLcBNYaBdMszt6xD5QTnem2exESUVSNB9LFdHnp6YXAQfm5wQ9k+E1aAje770hCto
5jKMa/svuSiJKz2YEh1BCNL6Z1nxlEmSeqimg+dfTuDCuWTkUfNtDjB4/Ody5SllsFps4bW/HmJ0
X89bMmqtb3I7FzDSay9f+dt0XHxlimFQ4aSD0pJjpCL2tAnhaKwpLifAHbXsbAntqCq9PWohhqNw
6JgIrlc0q0sRlWz91mHJXzwTC5DoQMYjyPGelDtpr0RjuG3PyQRTQ3ViqZ4JWc25mCyz+fNVreba
kg5TtOmWSqbvLojUU5Na+hUPYrssdAubEIhJHHBp6p1QxOIgioJnV18dD3Wc6arg4Xdr+T/2tORw
Uk23ie3fSIDjlVSzBcRjqA2cFmxhq53B0gInD6gaStjIOZ8btbJRgkDcN6oKYnPIhenZMQ5jW1pC
e27wyenTU15wP6alu2wxmgTsEGKDO9GFYjoQF57jPXpxeeI4IJzVlYzQf/UTXuohwMx1tpdSW/3b
3IRRZnwrrO0qWSrN0cmlY3WSgE6zAaS5fMcz5CemI1uILhA8Q05bQnmtsgiNm2KpT37C1EOpGYjw
vcRqqwHxmXOUjV0IIhmm4J2wq9VYKmSdWNiamxNcYugtiicsks7I/rvVPU44MOeY6oofimQN9qcR
H9IXMchaV22+nlBah30egjPwRWBUWrlw7K1dFp91LgqyaKCRnGZRLI+ye575kML3/wHAdwdXpUxQ
0zRviYUWTpvlmYcZIpKhzBuqFFFz5Cvh4J+4s6z+MvdGJgC1uBe8cr5IR7UOl+BJzYAZmuUiTQUP
EhNmRSTRMlZloFztrthWZfktlpWzr9wXSe2eygF5G6A0CMooGbt/eaWBXpy/AIdlczeos8a1whN4
NGoTZxNBNrra51xKchHd8+Zyhm1Y8BHUTIojRxRZ7s6/M9/vYc657lnvkz65RfoRkkRYbqDL4zV+
11WZc93HWNeDvJHvI1ICFXRkoyDMP2HxOeuvP/diTDRZaz78eOZhS5bK5hFfx2q1ogdSdN2ejlaE
ejzGKGnnlU4tM4rTcaR8WrwmNpkUFzV6DorEON0qTq/kb0bMk7/lKeiAG0Eke7Q+K3ren3DySQrN
ajP2TQzxYf2Tb8SaSAa1WWolFge0CrGykOFIxT2DTRL6KfSIw7i1Z8c/8BZzjNYk/FJdxLkFnRzz
WUxBf8WEbIst8ybAhyx45FdW7DqU23URBXAPPktUcuj5w7zcrgGZH12avPGJVNbQG2qwW1o0gwBb
UEwG5M0FOq00GU03HnialOoWEehbuijZXEiOQWhgBAjBuoLQuZECG2PV/Wt0wQ+zlvGCFwRBKWbM
rBPedng+g1DhAkFYdsQ2lY0UcpiYwvm2OYjVKBYOVxM1/CTpG5/DIYHmAd6EMptuuAMlwmhBdhyI
yB8go4HxfEXiQOztav4ea0dHlyTphLIFwPf7KOCQLmDIA2sMURjL+OAOl7MJPV7eoNq8960NbLcB
47l7ZewnN++acs0fi2JNKjmbWMBHcJbECjrKqnKCg04SUh5BkXIOrMMijXOJR8kfJgefwi/FUrgu
pSjwaVJQ8T/Dv3S1Lu//zVPIz0yDRoAEiIVldrDK8KfqsCO/hW2pEpt/0yocOsGFz4DFM5b7+O3Y
mTbTyGU5+fA60LIe1w0q6qs5nWsdiP3MLc0pltpeA7+t+2x3jBuGNX+dr8uh4WAAojKvAQCgJHgS
06LQvtacRk1GsmglEhSbPrb+XvPiY3hfxsQclpoWhNQRgzfrW3SEq4f7219XOCoWd9ygxjpVJzyG
W4+r/3jgNhrbW1M0nIgKbl6R9qciC/Qqmd1JW8Vf+A/zMPKnEsquESNbsrbz3AhYW02xjF1mpA0a
UOvYm41gQE9NJ8X61jKGXopaZoqOScBPY3p29lZ/jcyLeZFofpSCjnm3jqDJhIqWcXSo7eiOtZTD
Q9tHkKjZGngiaH+GL8r9qoi89F1WRsmkWIpGo4B0GrT2Ue434pl3S6ZVLcRe8iSpO8U4FTUC3wZp
7hZ8dVxECvtgW4pmMNub85sv4Wf+oYYnIuMv21bxUlblZsnvReunCuh1TUKN+/mv/DfWyycwT+8e
mzgeNGbdjSEtRhe/MHh8sE0/FxsTouFqDBUQHuaygdFIzZj+TzMiIFjd0XDHucgOF4qUuTCaiRZj
VB1W8GSeiO7PqFia74qMrjGkNB3klO1Mda1nLWXBODCFtKv2sm2WtRIpqgx2cs4GexxOGU1ZjqSJ
pgC9+Fx7lqEEXMVTrqJcdsgRcVkbBhTZAf/vIj4DALwyDr5QoJ+3dqp/0mJWGnRq68Al53/6cDtY
uAeeNBbGqElbRkfkoHFQI9T6hg56wAu4Aix04x5atGdrn74Pqf0F2GePgO3hQ/gDKlDINlikxRUz
CwXPquvVwSqrlkyB5oyFrfl9vHymlWNoizJ1hB23aFsa0nYOUXraqZ5fN3vjkyQHsfBpkI1RH/rv
3rdM2U67iscG2xKAJlwX7x/AJMUD3IHN/wwj8UAuwifSmw3rMSQExTcyxE4b2Rlje8VXaGiVNp+z
QaaAIRnR6iXMEsD4U7zhpOrw6Y14/unrGSscpHTissTHiT15K6QsDAi6NsUuniTzLsUt2kYLADCu
n4TsKSsLNb3hyV7i9dU2fQ1AgREuvbVbKt8D28mT1QDHOJRDk2rxZx9QKswTOrk3c1UXa34ZqJwy
4e5NtmPw3QzFL9//LQKhOD+ph/pKbCSiSdmvbynMHkvQEvR4CKZ9cFfizLmjG+CnXv+t3J+xw24j
DxBlVl7WLo76jSOpAJwrohP/25jtjdEj3923iMQ4mPdyhlCbCHBUbf0FZeUE6KV+C+mjGFuv+x19
zGbdRiC0NPo9dddMGHPfjTXCQFLkBn3AFjE8rp3Y/C+Mk2aNAHp68qfqpHWaD29/h3zGoxY24Ytm
k3DYv8rFKd/+OxWuJgm/PBeMPmestI5YzCFO9QY1uwvKY+zQniyMe5lnniQ9qJTvbwrCmuJaxtCo
qtylc6JZBncG/xX9QdfYuF8Q8uitMrEZ3TdaRyfxUgoRUMxGUh9c0rBUzTzrmFNxx08/NgCd5bPR
8b05UVTMl0jP4za/iwrquo9YyuzqTCoAKT1zYjUvL22Y0yvSW5aSDng0x9xwyCuSiAuGhieBKgPU
GKnPmlxg+kF60kROsLElb3COe4pd/QB0PnakQ/cti+91VgCIVESdhsFMr8OtEppCkphyJETKv2Au
zjk6ghgYLApaA2PCcTYvFepqoXwl7xEAz0FPRVI7ikLSllJd1Sy9rMUZU2s2rtpgzKY3DaDYeB3A
UjSlShmDbwcd2HoQgiNPHazAePvp8YiuTn/5x26Rj6A8YdLjKBk9uOpzI1NJiUhYAgCNHYgDeIur
DnjCsF2yfH8AGaWSF9YBHGLfhNVOg4tofHtSerh0ZRO1bHAuhVBRcVel1hpERO6GVUiS4FA6POD9
vZYnb5/ZLbqC0vNixIqz/lTR3ccxIrve4jRMmzLgD6UOWcDdTsJUqRTaruW9Hr95+AIUfYpzFFfH
caeN54lVlNOKWLMrZdSZzmVl+LdAoLBajIrTpGHfLY0Xg5ZGwUsJhGoEjphWVto/fSCBkfHWfLo7
kWa/spPPv3zTM1Bg37xbefDtu1f2qxe0U+Hnulk3ry6p8ANvlKtpDrt7/1wyKnFClJyweg+riuuK
c6XxjEzzDS0vkNxDgdSycIshOUP65TBNavOnJN9vrODKsX568Da/SrsmvFaQjLMqN70e7JmYX8T7
juw1zcGjvdts5a5VuTDNLuKLCmG1Y8tOaIASzEFn+HQ6a1poWgIFBuz6/Gl6YSy1TpSiAsVnTDNS
bCdiTAtdq7fY+PBgDpba0xEUAeyWi199+U+1Ssr91xN/4RbfkBFQhqDwXkKr8faZxJombR9m8OUN
LOTdD6BN6tulDM9umMXzbOV5WcYsyFV7AJX7tZe/UfBZxLb9W8nQ04yS0Co1miZ15yVUaT/VLzPn
AUQgoBVOvLschnzBaqDQWXZcVpjg0G55/9Z5826YEoJkHOgRavfs4PxluLyBr088rDmP20z+6Ucx
TKSrlbNj/Igzth7mOFoYCy9O3SOVgWAPcQFwTF2PnpXl6wnThHxkBh9JNy5aQIxvs0O7pA7829Mm
sBFhj2zVvDBQ0jJKyk042xUo7KbxWgNBVq60exPPmND3MNIlo2dN21OHK2FYWQ0pjoOxjgiNZcSz
she1mA5808606Gr56EC9fif6uhoRtFypuskuiBcyxwaEW1PZTwL/VjXwLz0KaXOik8qAOoCD4HFC
ox6HFUPa4nO4PXOynNMGgSexkUYcuiT9VzQ8tglV26gYTGAoZE5kbc2TTft3h7exUuYmOoUCUgpf
ogd83IPQHz+b8+x4f9zA4Bh09FopXTPGrGwz/JocwqgHDvK5qb0aRFfZM9cK5AW0k2RaJGQFjWW6
Pn12Dcc3JLJyiy0kcwfwS8himL/4/pNs0LCeS2Q5k8tmumscy1I1xq9mNiTkm2DA/j8DxqyZ4z6O
SSp0DVH/M9onRV7rL7ZWGljJ8XUz2jDnHd+uzyORghhP3ue0OZaPnShqSRw5FESXSY2tId41NHEA
c1vMxATV9xOgxtLVhc4UK3YO8mjXo/j8ibBzB2wZnP/isicXEQIaP7gOPlB/GgI8kedBSrui07IM
K1xYL64pYk16bi7IUcG5gKMAaQfzyRlgghXckFilETpVKhOa/Gut1iajVwUm0NXsTTFPRVB9uyZL
zcq9zl8XfgAdmp9KGBQ1Youd3c9nkZ5a9UYV2Xrvln5mMEAOMopXiG7H/eVmwHskuzm96ZI5oqgP
oCzU3dNKQZhSMoO8SfEA0G2oaDD41Z9j14D8BqKgUoSZpZpy646I6iHr+AFAqOxpyil5DFLJ8+YM
in0Yzl7ShIz+IokElKKIZspbf9LkVGHGnoA/XbNPE7sRAiZrbCSpbGf3XVaqcmTJdiCTg1BggTCp
JLdwZ6GI9Ux42hAwjRruzqDwgb0wIauivixANjPd3y7HpPRlXuWu+yEUBsdYw1EiC12NWDMAB5Ta
6EjM/D6jLYJrqoPDd1n1ZZ42bu8bC1brj2V3Tn+zDeUgUGSOmEvWYyIBglsCQlnG6+EwXXhU0aP5
q/pa9bOXxROAxy+EA2DLjTm09fDd/MGTbxb//UdzCn2Y/EYIZ4o1Q5Ng7tbU7sXkxY5JmEQUtH68
TLQVVSSyHPcnYN7NnKyNjBdaQ9VhnhsCJ7/nKHPJT3AaHBdgId5e0HkpnsrEazgLnBRsVI08Um+x
m4jAyhBpaFfJfQsPGCMonbS1hk43JIoe+a2lnVoNnG+MFUeZ2I3rie5GR9Y5GUq0xlPMxUn+krg6
Rbi5AloLw4ymVXoWBX6JMW/6+DccldzWotxe3HcyNDgqHEi7T3Cb6i+jd/j0kseoRSYeOsWDpCdb
XtN8UE+njJS5SnwqYmJvj08edki6cvYavcqRrC5G4XexPuUVkniVb1z/ysr2j/rDtem+woAFMvDe
R088/NwCyK0e86DzBei/ktYrGaymqdJeiteaTifSyCMwuehP1xv3FQJPx7AscbHf/ibdZmywKaW9
ixA/cQEeUDxp5egAuKz7oaWW1MiNeWhJdH8uLFvoY7kL0Qdz+0VFyPpgdqBlUZYcZcABkMn15VQi
NDwayaMBa6L7EXFPkR80KAa0/e/cBKKmXym7AmhVHQiG2FUt2nsjv8FHNcNsCl1teKje441xaAEX
E/YrfL+6jpnksNBdqe1hKiBcc6rHAai06JYTjrZzU4tAFvS70Lmr1Rf6cRx0mGlm9d8C3xEjtx16
q/lX8LlwlFL2rqVNO7FTRyQ14cRVY9+kKhdxE8+GNYqI3poJ/TWOFU2yG2VlnaFDm2go5lfYGB7D
JABIQwiLPB9UxReDxlBs6vuu9g7yNLC5XNJStRwUCFu6Tq0HnL5QLEZYubv5IhAPLAJAoVtatjHH
FMnYIc4gOemT7INyIS6l/c5Oxv0PotIX9/XAJO5G6KynsZ507wwW+goFvp5YN+nFm1qC3zuY/nc8
lzZZ4LDpHI74+1u0wUSnM3ZfPC9TTWOxiKKxhrEx3+YYGgBHRbsMip35satcYoFai1xR4GNozRiX
jTMYaQrKTdTV2/2J4S6ELh7Awww9fFS5lBczW2pULoGI9RR09MAR2T/2gbLRN2Pf0szpp15NAypg
8q+AwB5M8QmGJPZ8OGEQwiUdREGwXHq8zgbNxQJ140AK9rURQNVNfLHSIPYfEHv63VyatFGdGgPg
Sc4t5ro4qVJ15rPBT1TsMyFCOk8ssYoO8wmTRl8GLWXWxdqU8DeecsiankYcW9lV47iwAWefXbAH
S/vchRdeA0H2e+8HqTwYByltptwq2kQ+NJC4kP0srlG9w+eMJNO3QTZxIEqA/1VUFw0SnoWjSyLu
kk6LXF3rps7BE8t0jQGZZqK5vCehzoKjO1AukhUn8tLyVyqoxKgrw4DEQlJZI9PkPL38Y/51oNFr
zXIImXgGA55M6y1bcfroOq7htq5iE50qmnd8AKTmZ/TeA8Uf7Wp/FxdzwHJKwLVAy/6EBBxv7Xgo
YOZg34cC3A4ZCpCUI1k2MBH+JHzn8PgmwZgZ2grCa8+/p2zILNP1bORDNljzvz65kIL92U6bFdlN
8e3ejSvhFde16nDZXAZ/tSv/gnnzm2l3I6OpW1b/ySbS2gfTN8OxgpgfdQmwG09PmCQwWuetQe6s
wveQGn4Z4shvyPvtUzguFi7kWKAubm79cTKYPCtRtc8QYHtoKO2UcP6C44wiI6x4v3FVxGS6Jivs
DIWCjLw1yIVFzJfo8RP5SJ8S3C9ynfMjrbG7x3SMO5yz1j7aFT8+hzIVn74sdWgZjd8GiOuJp9+x
Js7ghDrCQMDX8uYCKnmoyOSeVkBHAQIc0wGdZ2DaIv+5rUrvp4Jny+Iu+DAq6SkEgFkuavs7UMb6
3gNDQRZXAIoOWdt5BzhN9mjclSrIwueuarh2L0OzoeyuFcCGrBYpQjcW3WHkMwJlRZcNvl840Hiu
MEAx+4wQPRM/1YzyUJiul+Nd5wZKs4eDxSmdO/iKBlvMh66pN69URnXIV/Y9LtjHVhypXTjU3ync
MKs8A0Xt3vZednzqdehrvyh24Ngsbfc7xzAhqiBXK4SB0g3C4aDO63q1i7z0193w5pC5rR2P0vTl
TEY9ioD3X8T2EfJYXwpeTZ8JnqqmQnzB04oTgzaa8wjXTry1e2qll7kHFXNg8WOFUjJSkbdVrlEC
LiZNTeyLQRei9Xjb46v3qgkoDk9q67/v/yMOMrjO8EqzQRwPUXLYVlqMaV0VL3DNVcElOvamSWTy
MzMa3kBOjTWTJQ9a5MO5UxK9OjG7fNuWihesUmGCdyPlGOPk2ntUihMI7AWISC0SyOkq9hRnhnt6
4dFfQWffVz1Cjhr+so8/MXKuOV58gkrHdeX3LvoPEO09vQpnLsdLha1/nHrarCOVaEo53ljOWVR8
GW9aviU83FynrFGNmXPTpmtoZo7aXr4u8L3k/hKs4GmEJdcwhNCcEhbz98Lb6Mg8/OHERpgk0w/o
xhZdLiTgI0HkIjPIB6bpNYMJGmpuyeRAwhZ61Xrl9gYBjfvHWXAUvgJL85gOBI30TI+UHfRBlVlQ
f6Knq/VWWUE1W+mUn5Ax5dXTDG17AHvmCTAgejAvtpRwK/Gy8CZv/vLgFiilSCX0y8kOtWUnNquf
UQRE+FL/dzDB6oJ1UyRPA+f3VN/2oxPvYoP4VMBffUtK0B4U/piooihQvXDpBFnWZI7LKaZz4vBC
P9ot5WqvnFNltJCsq3Q9t1U+g5vd5WiBxLq6Mu6ML1llr+dxOxrKY6ByaAuJEor4MSH7XPZQj1S3
yPWFQgf7AakRs+kGON+bNcZxBgSBGVBb2RThWdZ7O60fbzamL6SVHPSMT2nvcpBVLjxqmTn9j7DU
K/AHiUm7HFjiOsDXxLQdt552gdGwJAIMQdw6SXfQtNIBKRryTI9g289Q9xjB8BroGFUQyN57Y2nA
MWGk5ql7LPCcQrNE5T/VQQoz/xX8PBSanJ39hcLFpnwfljYxhkMEFr9fr28EWPTIYLZxK8LTeM5V
tiLqFpDZPbNYDvyDzA4tOpkoWMx2w4gY4UGQGoeqb+56WYHYegIfd6hHYWOUxbXosuYytuhfNmRI
Osw1jAeWpv7bl5POAONdcERoMa3mXuNkfAtVXuHe5MExzRBhjlv3dx+8QbWqE+tBSaxUhKb+8KD8
qSgRxlAVSCQb4t3ATZVn0Fc+5ooaC24QaTHjQ6NH1Pc8gDtEUP2lwtR4NlOVpbQCTJ1y0+mc+5on
rMvN6YlwxEHplzHPtKf/lUvJoGDPIIsBcldllO2ZJVcqjlYQH3G9SyBhr1Ygx7SnF0B/NXkga2IH
04SzfT3v7dDNqyInzseNJbFEL09uYmMUxEIFHfd+HRf1J2gZ3p2Q2tivcQ2udUgPyNlCvdXdKYoU
51+dPpfiIpc2d/JkCuifWmhQHbrUw8xr07KArxjDVpWAJHSUYnf/gch3z+2JbDu0+zEjRiaMT6Mg
qWUoNMlmjMRO2OpcbQrcZeeJiKto2hzMfV5AyeowX9plWceA2Y/FrFgeQnRSI7zJfvT8v+tLa59u
VSxdBi614agAPASYNqEvy0qcL6+88iOUqZntnK+ctXYYE4AdEdm5x7BqzaqpsrhkZNCm5Hu4sIkQ
cX1zIsu8Xnc7qkXTabofW1LoBPF4fboCphq0e8cGJtfxKF9W/ff2GqLitdNzP/ydj90NXQ3e2j4o
AUT1+ZN5eBzOMUGYer2CHNOprUyg0FzA+PpYVyHDqkgZw20JizRY/NUinsr5T4cc5ihN/8H1KGk4
Xl/R1PNcIJbcNGmvgyV8eJ7ziIYyqdBIY/Ac49ob45ObKyYRPNUqJp5xKUcLosSDU1Mg5NzXq61P
KpivC2V0FLYp7JpRwZce2sWlHjv/qEVowMUGaCfFiCQXD4iwUwd6sprfanaY+bDmXLRvq948qbqz
ZITNgmq3dlQE2anXFgooMpKHdheS+C+a6c1SJK7fbtB5HaF3RkOqbiJ4ZZo54Beua1ECQzVSYMNp
wI9i1gN0OLBp6X+j6NzNL9SgdFoU1za3CeLsbhWYutkyFLxzUOKk8dGAkgNYnUla6YRQiaau8T9l
//6ULaGJ/m8m0kSIvaFZnA0mN12rZPTYlGt9dFy/839HO6cG9+Qhh51zipO0R/+A5MlgRqdqpAW5
jketShkx7WwaKHt+malFFUbsh7dz/iekEkQjM9ewqO4M/GE6DtBCTY2IukKN2CbNFIWOkUwMmmmO
p7PJTCw2/aPQjkMSTesYynxhI+feX62pov+RKjZFRlWhvvcq1mUlFfkrhtQJEwUJx8cNyTVoFYWd
lRttKvfzx9hwooBo5dVkYTF+4fygBtWPKETuXSa819XnbHwgrljVGoauQlrQ5/uyXzXE332UtdaF
lPjdytdFohZUnjOkiPOU4lD72CJjKAdVn0mjDiLHzeJhnfLZgDKSGvmBTePpKYeLOGiMtDvm3j3b
Gr0HnIto19hHP0Hih1MesNguQneKR//m1tBJ3/ad2L1lTmGR9o2ihmavc7fQZQkgGyyNGIXbCF31
bFIiPMgioU1xPxsGST/6eKW8ow/PoBh117LgRkCvtg4AhAA2DbebiPImBzCw79uubBUOKd8cX9nt
oZo9fnoEySGtV61HjrzwhgBe4aJgZiur47xi/KwoJcaYQDAkg8DLRfnQaZNYpaxkER2/SQwAExze
JhPymQLbfslBzUcHLE2jN0h8FcjYzwhdPNNtRBpX/+AOeyjpbNiN1/2rsDTC1NXjx4qjwn8LfgaI
ooRRGG70F7LGIT1jQg5YZmJwFVIfinute6ez6OYH6QkeGDXRsS0gwxThIezxksmS/lw7pTKcw32R
ihpgDFgKhz+i66PoiGHAr5A1J2WWzCwgcSGQtO9frpJQnnvNsYDXmcBqROfTgXxd+1R9kdIVCTpj
L+Jp4WuuF+W2XKUSAHYMgkKWdqpNw3GUHAD0VBb8YeIAgM43OqzwRt6GhOzxii1airFRIRFC0PVL
O7RjsHK44MstPM7hogkTi4eTHxXrCOI9cFO1MoYSBixXAIPny7L7L9356OsBqGaAix8Gh3j9lbg0
/gejWwPG4x/wIVAQ/j5mv3c18abO7KKdYCuNbhTTHRT6wVzp8sIgIcBEOLz+FFQkMGN4Owrh/mN8
mNYSCQ6M/T5611ayPF6DrLMozI+aGW57u9xHnhFkpuZwmDi5i/fdOrKtjAdSKoeslMFsD4yFYHzq
WVRMJ4FwbFhysxjTFIHJ04TFCs4MkCj16WhtVx6yCslpmDllJwtS/ISy0Rhf310zdHapWgWEgvCk
Kwrzc8cixP0/FDIN+3I+uvVI8+P6wRMCx1QowZ3Y0tf9N8ZL4W39m+vUB5iKAECP1I1IN/hNYiaR
TXSdDtpyk/1V/bpDyhfguSCgrpfJXuzsCePKGX2dIyCKVLehOZy3b9bhnvsonoOnvfpiL8+L4xP1
jStXXce50io0j3vjzhS0bMKTu6XiRbXHB0vDa1AF8d6xQepdcE62gqZfPdjsJBFzJmYNAMFgc9i3
IO2wGTMDaXVNfIByIe4Hiq6qhgGLL596yni/o/Q1oZPdx6jGAmDP6i7d9Ld7d/3etQLcN9XAjSld
uDJfUdh/lwrF9vqdIoTaTrljMf+U8oCT4ksFA6Y04sJM96rXT6Dw8QS790BXgif/HHZghE5l78rt
tBMVaKaIVxCCHffO2jkKsJ8EL0Xfi+dkQ/xjzM1vCY+eDycOjaljvy+whmLccoaUZfvndMeh1U1d
qMuhpnaPE+RjBEaew8WwFkq8SQlSUwdHei75wG30ZYRuxfKK07l1CoP3WVTqkR4pnjjLKhDQqmET
NBWkzHHN09qAbqrpUclvCCzTsWjDu4i+SmDGAbl7rF/cgJabTVE0d4/2y6ej5Nrxv3gkF3HXUFfE
q8qrQVHN13D4BXkftlx23osGLbxE/z0n9H4HW+PG2w94+Rh2rZVtwcfb2ZYOCd0B09o09vz14zP0
yN6LsHPbfkqaLxxh+fXkOFbsJ94lQ0OieYLx4CxZ3zg2wxR/H0kom10YyuAOZJi6/pe+T6iqvMI7
DO4X03LEW4SbxRCKsNfmWg3OKuaNdUM5jhp8hedAiV7zEsxOx9B4QZvI2wkFvBjEJ4hllZOMWtDo
djry0XaM02G49JT8q5RkFQN0kUJwquz8RRAmfu5XUCfi93Ut55o0xBzyqZI2Grixe7hu2LnGIXRH
E7C0t8/qSKUTtGngIEkT+2qu8Lj2RBU8n0AHr/fn+nkLRpgOBTJrwoGqOU5wf255sqYt++XVhgwG
C23upQ64N6iMswGZvoi1zPC4eFJ0vz5GlgrNP3EUffiE2uYKlUG5y5mG6QuDsQKEYZaLbRsbfgzN
8PE3RKxKRnSxejt/MM+HWIDs/dV2Ooh+rwNz8TBdyiUEVuk9+dI+RyTw7anp/FnNOkGYxTftMy0x
EfNfXEU1ghip2DP7vRu9HiXCwj1cMODJW6iLf3zBMNDWKcH4qwGErt4gaYHramnL9g8UYya3n0hJ
ugZsBl8+GI03hIS2gtKk6v5wXgrDJ8KxZfK1UrF4SM843h198Uys1O4j3E7SyvVJugLRscb24VJm
03rhhVEGDOa9aBLJnvIY97Wi0oBbDlXTakJH9TA9w4wzin/6BS3vE/axtR8NF9uuZczNmhODNDap
A2PwfDEjliCXOt0A/ehosc3nCfGiQNFciWgxY6S6WY9BaW7CzLcfHF6JNjtQM4XiQZk4orVBLhay
0lWS7vnAWtamACquvIP42srE05vSrXzRwgAZnzybeiJ2ijUUU5P/IGXg9B1y43KbtqykJXAr20hv
slg6fkKppzg06HuSJJXVHpHLovfkywmVeJWsPsO5EmY7tgwFLWE3zDL6DLVPvRN1cr9jhFy/68oZ
qwJPURz6/TboLRK08zpl7V3QXfKaPpmf4mNL5ND+NbwOmSyK8twOSHcCz6ZGbcAZGFdWPQqCHSwD
IGqCV89t06wDDv/dgqKzFsI+BA9uB7U0oyIRBwb73pi/mz4bw4Zk4C8yQGSH78LCNHtrZPGurZ8t
+5GxIRPBc+vT3aMrJh1nXnGTNPkkjE1l5Z38F0jTSiDai7WHFhHE9nI7v/7M6gfffgAsnlcBVEZS
D3Wv7jSyfqsb/zUnKJBTeN6HyDAYtxPOeoP1GK04chqGvP2514VOyCYbX+3fQslfb/TVMpji7/n6
porbxyuuByAUI1P+mOziBR7T5OCzHMEFeN85iefCoypbpwnwfniGZUVLKRYUnpJam2Sw2EhInVCQ
mYcNjy61XUDd9GAehAzAkQLWtp6kgmGSPbEKMdzcZo99nk63DE5VH5pj6MTcN9Xv7Hn5t+rbQb/E
n9F+4k84LwNbSheGsVLDHirH2sIW+tNWZmbpkoXmJJvrq3Q0IwUNYjdhJdQTj3m0CAa9+tj3hXA0
SJ/ZAela+ZzrIDuSqFUq2hLz0H5s5+tGxU3ehK0GHIWnp7PzahyRFNLGgqbzu/y35mda6LveHUNg
UP4b+3YMRPnH4zUXJS62TlnPSEr5xY0Pg7h/BVAL6/P+u085nRZOPgZbPPW6r6hL56upplkQE5Ja
fXvOuiGTcJ04yvdn3sqj6kdUo4utpbWznjSGTqbfzDqcwMx2M9mF8JV1wINiAGCNGESCNCH894E2
bcK63vqwZnDqrtOYK5zHiu2CIisdBKPjr4cALAOZcM7nKYlimoKTORsm2291vcZ+0bPxUO8S5dcX
ohPIJVCn64TxFY7btRVm4djomDiFQtIbR6usQ+Ichel115dOo6IzT5eRm0vwieFaVYIfFjhel+il
X4fZ4CLb4Ub5XquZk8eNiECgEZu1DYg3a45MR+bCmi/uOsqAHuTjSc4HkrhFB4d93DfMjhSnWHb4
znoVlSdOhhNMl5tYLTDgFRwR5FOMsVdi1fOq8CWS+KQHc60/+XRiLt3AFvBQRoWWmX0LNcIqjIBs
j1bGtNrbsM35y0yFwOzT5wE0Wkgf3+kDaa7F2ijdr71d4S8z7wEPCd/iqFYKOiWr+AiOADBWVDC4
OaWotm6S1yBY80PBLZmLi2GPtJQFbNbfDMVp/T3TlqvRK8orScaPxZ9cVhqPTk+/5HdeJQCpaeHl
asB/F6CvONArueIm+T0WVHYENu2VtHvgK8dR9NBTmveQUSwt04eTfET6t/9OBG1BKSRn3pnX1coh
GgUXVknvVsZu0FQcdKTOaTVimR3IoXrc9wXyr7QeMze91CyLQgFaiLbAxt5o+0FWd/3arsa4CfmU
Bys9ZP+mC8ZsuUzjQ+6zqKQ1W6qwzq93T1mQyim4rcTMlRBtPDBtTZWP55qVmgMy82GP7rTspJWK
JvqvN4cXmWBEnEdWVSfwO+zS+vv/Yjl+XsPQH9285q4KwKe0fIE0HFxO21oSgDUh2SYwCycYTkUR
ehb4B0qGYl1YmLnkxchwRJdHR4xm8BTB9h4nLaKuuswtjxd1kiORU/fN+Y5LOUGgOq+kQLLqSj/G
Z3oDOSHlTfO8Xgin0Bf2c3qL7LCyY8RseGEf5jDMw2b6U1wDVap9Xe1V4BzWsxqIjpp0ORiM+eoY
LrcpthW7cIXcuuYUqzmgBpjpiy/N9aqnOQEcKcO32KHQHUYyJz5jRzLDrNEYmJKSKWHKtRf+4zOF
fNaBFkfviUoFZ4kcevtEt0XrZQ2L9D9frKw5/bK1mTTatvvIuoBqPMiIBp8Ppgza581xxZDybirW
PU/eoduHPbk4cwUWdfqD3mYQNjza8Rwo0NoPn6x6w6W3b/NU83mvYRVv6PQzjP3MVxASBxP997ng
EODElbfmbPFWnqUDT/fWKXjS9Kb45c//CLLkYtew1j9+OlWdBbkA1Q8veUM23le/Ys9p2/O6/qyU
DaNhiWsEHPeBfPQEopsnuK9cm8uw1d4YpoxIh4y6eIrLNh+yF1f92vvv2Vfenn287t45kxa2bl7k
7S14ljmQS4bPhBL6db2Vq4F2G4hCI9C9JVvANshtgbp+h5XLEhvQdktlJ8kCMorSoVxcTJLDHkp5
4iShMXNMIYybmbrMCPC9hSpI5zMfnGYLhUh40y9FZS0Lhv6Em8VbyrXmNUrrbcQC2pQdvEe+cjlZ
1iBcPBuuP75TdKT3ZETyPNIE/wT8QSTf7IQcMtCUye1RvO/W0VjlLu+N/s24JXjm24wHffiScAfG
we3jWg+4g3RV6M7H+h0FZN58qf1pRNlRr6qaip+8bJL3bq5wJO+ekW4lCmkQHJPnKzgsd7PwG+v9
bFDXry5GfKdJ8RK5QMKA6c9Zuppyqf/dmKfgfZRh24hMlT0wIZWqYWtGVh4MauPGL36UPqYKBqib
+v5H+vM4b/Yt0rwrETgYoWpXZEhkGfnXkx4ZGXH8ldse/dZJyUB0UT/tHZIY9iZwT/3WDt8vfiUR
ED223KLc7PLeZgM0tOHJoopvadeVjfRHCjHUwUZjeKYdBhnna1C9jcTy7Y4UgjoBAV/+SgNuzuML
x8WfFOqLnejz4FVkFT71HdpH8tQdRLn906nYw6q2h37LJQo2UcXcfE9hdzW7VbkvHFra3Lj98ZQd
L+BewAGIIdvkwUluzSPxXnQQvv114CFopjJ2gCNS8jj89+t4+KPWyvPiaZzhE/SAG3ys1BBRWG8X
WySKtCjHpbwnxAZjdhR4sJdRQx79vBPGiIhj1PJ4vIA2VsZEEtYcX7ckpBNbBB92PvDuuYGV+UkN
gcbDZ/qNWhfXUt7Q8rnU8mTODnS0KrzR/j+ZFYoULlU/L5NVbkULWu0nlr2C9FRcRCJYQx4yMaSV
Pd3jBrv2AymWJ2MbQhlg9ShxYAXvxzei+Txcz/YlBUMvb6KBF54TdUen9ACFo8TWDuISgOxOJrSA
Lef3G5zZrrjrO5V//7c9cRlQ0836tkWM67USbIfwORzphYYe2nCIORs5+f87E+HdbqkHTkvyZW5B
z3rWMP72qwFLktELvvZBnPe72M4QyCNKt5xQEMKOlB7j1FZAhiDJVDH4ClCRozzZZGphzDF2BOmu
YWy/hBzTw7Wz6GUNsiEMsri0TEU5sMM79TJbQWBIyTfpiSYVs8oJ4cmYi7UlGwWkqWw9o9451RH7
eJmwrxkljic5pkJN6XRM7JzBHLwZfLc/oQ576RwYhJW9u1CcxTZYtp7tiWtJ6fscdsGKL6LtoAkU
4VXR9ELNx7W4+B8fm9bC6FrDk+q82aQOBVEPfamvclOYG9dadGS4wYlMd+UycPbM6ffCRKwGqaso
SoBOfV7xr3rCEMuckSBwztQAjqzGH5NJU4j49RzuzbXRXXDL+vN92q+1evFNMv8VYeqQSMK+3Ioj
jX6erG+m8+gaSdwa+FOkwv9KKoiY3pru5IqIxr1PuGxQzPg/y5WzxbifDb09U/Hc7J01kj7GgSf5
XXrts61GTW/SKbxe8ElNds0KMr/lPDFudTXbus0vynSFu46vfCUGl1PdWf8ENabml1qnkPc6A3he
wrrrEDgAxwOQA6xYW3Vbu++i3hyp+rJgGAYbaa/dKki6GdiltH8YcLkditJY6yfiRnHr9DIW/z1b
EkrCdiUmE94KvdW7JM2Z71r7qhJ1Gs/w3XOuBSKxCL+3KgXOY3erL1Mt21eHDLf3TC8wRhiF6fT6
oEgP0zp9LtXKEKWOEM4uH85LMX6nKAdcbbJjRiHT6upYiy4b2x7hlQGjfGBQAm4RNDfzefq1A4Om
EGCmVPSXEbeak+/B9MxrbpSVswYstDxX6P+rr8y9eTX7c40+icbsvJZj6GCglh523hFsjIU9xuk7
ASVRAbRpQTODlrdG1xh2gQoflbRBQ+DDkKA5P6wS7r2huGc7BOnClH/VJutQeT8WLZifxG3NafgU
XqgUCXYoDTbeWKZU00UvsmszkkUX2ocmxajWGox0RyoCGLXpEwWC3tx4wqWxTZLn4jzbKpxpkVcg
CCIdMeRT7FqnYybIz1X/KenuK4AWrniGzE3HVhH0xl/jdC9T2IVCdyL3ustl0/BOFs9xI98zUFDP
/fc9JPsBRyQll2gRWlOKtVTpL7uWIWHmHEOz++TH/XI3dTpAZYJe1fmlGtKYm4ctTpW9uP1cdOtZ
6jvwaqrzSJiooA0hBzLyZiYqcmCRFm/8PFLkae6tZhaDuhrVIz0gEistpHumjBMSy55Hbq+D0ANt
D87hWpswtsy+H/uL5N+NNKrRAqHU8AKLoYP5GjN1bdQd6EnN+Rtr1sDhNR4xo70fLxKUjSSiijbH
7c0btSXhHwmYohMFxaAX2AwP0S4xt3Mi980f3a3Fjv9JIwy/o8movaDGYIZOMo6olR3M6iKuPNqR
jCf+CZeEnxFGQ7040ONayy2mw3tut2Ncmu+G2xIuDCIZXgWB4fgXodwBmg+dJMHvyAEb9P714el7
0OJtxRMjf5c9SiVlFE0CY8AR7Tan1pDdtwysArpcpeA99CfREMXV0WGXvqyTrCJj6R2HYEqYFxyE
9zrfu+E7sp/MQrHEjoeQo1rMaA+hsWfxAEqDNb+XhPP9t4BwDq4xZ2FXxbY3EtIuaNeH4wUXpO0d
35GZ/SEFQLmxP/FmPKIw9C6bhJRjqqClG7+hF61KK/dT9m6AQVg5nrrSZOcNYTodQFZDcHPtwOPz
BN0nEPGZrV0Fr9fmih86+b+L1jWXZ++GKXNfzaK+BM9PJMUdxO5N8qV4zEqHZn3/udt3EpZ1Izku
BZRAL0WdLrjyzfV1trplwewHlofA5YjsrpBcPCs65sgBdHB9mBQXmbpNVDHTKwZVWMZH4fViC6uI
j2p/8aLXLUaKwLvIL/wtvasBvprhWOSC0woZ/KWReH/KMg7P1y93Fx7VfjNBzEn6snh1xB/0QS+a
EOMvboE3b0kIEglQqU2w8FbqY25E+lsxkO3UjvjfDPivcnpinSRVV7fnYMVj0pKLcHegXYPBsbaN
z3GnS60YLGP9oZrh3dFxVbAmN3VzHODthFh+vQTkFS+LF3tVg7EYfu71p/AN81Mbol1uxjTnLN+e
I9U0azVHOJrokiTnFXcuf3b6PD2HjnGzn7ZqI27eczviIOy2b96Vp3t5zgtwTDENm3CE0onYih7y
0bewwlXaPJTHdesCA4KhZLXg72Ww/7pSrodO1UxWkuUEzWP+qWPE5EoGzvybTwC0HrtP4MbAc9RC
2lb5LZYjBbcF2t9lP2TNyVaJ+yd07xYkBEwRhtoiHKc7ULDRXm20s9PJgM5/RdigMthl5r6N71eO
WycDUVZ5jsIK+ZgItitYWZxY2uHsMaoQQ8clZ3PZUOzd+WlvdH7ly2cFKk+vt9sfvHv5mfsZvVb/
w0sIAXeXf8xSgKQfnYHLwA5QIczbNjvZ/lZH76CN+N+0ONcWpjxbUS2oMtQF4982VxcX7PE5iIvj
NXKO7IRzaF5YC00MF9Dq/xZikwX2HPOcTYmvzrqI0/ZjsHX4r2LHox71d6t8znCZ9yjaki10C5dq
xNVDRuRHuibjt0fBmEd9x3vlud1S1ieIux4TysLAKaecTPph6NzIzpBwyQRUfsP2hw9UV5Xngrya
bOdrYQNnPeFHNq4/cb1LKnLUI9PENVI/B4k5pR29L5ZHcjqY9CXi/Pb+aEy+pX9sE/uBercm1ciY
pF4tXonlo/zC/uXLWgFYat08ywcL9KcCGe7/FGSRk2Bgp2Qb+QygM1ohfm5Pnqox9lIIVNZ8nWn2
7q4mg+FEwl2WfzRv04Uf+hXT2qWPrYeHfA5hPrikWOqXWszIvhP7uK80qes9+Y30YqMvvBcpDBxS
XJA4d8NX3is0Oyi6Jg3iDULx0JfdJ1Yw3pswSeUGMLq5GB6UYk6Pe6nLlfVyhe2cZFpCYtZ3Lp4F
wKc5SP+KgqcmT8YOVI868ZB79cBGRf1teRy0e8KFQ1nvoZ21SKf6MGX5023i+FvZ/3Mie3cqBvqg
05K+TqGrqCBUE2CBiCwCmew55Kl3lOH7HEcklMMv7VNXUuh+eG4R0BK1Ga7nK5d+SGnNGyJl6YEY
Dc8wqExL4t2mO4Vu3sN7ApzPHkXrI+uvCFK0jANDhh01gJGASV2Yq5FrHDjv7Zh2vWadl0tBNK+x
aJbXQ2MVaQgABwQzFKkRgFO7UgS5T1m7Va9gNl2eb8ox3tbKdA4BWrBHA/BaeaIV9l0sfMv59GKS
G1qL0d0LNbk52LRcW50INLPJUrCpif+LR27OEvTmr0XTKnRZgYYXu6TIEpTrCuT22fBZ/5jm7mcx
Aoh6NG0XKKO2d3wIobkq0eVpxAzigB0o5VTQxavlA4L/zV3EIIRv6wP930s7es2hWg+AveIhglQh
aZLPwlNwKNy+qkJ154bGF5ezRBpZMX5YtcNtckdBf5q3eL+hRnCrz3VyvIGO3RBNmQ7xJVsNACrG
Ju50Aon9mVy6FdIfCGHTcfZXYQ4RD08Nn3E5/g9D+A4BAokOh6ghHlDGQsBinyybYEAL4SgVwENh
lA8ttJCVevmf/01G4V+RzbAwasUFE9/7cyLshOxsgFY6g8ovIaFt6oPh0lFXu5rsnhOJG9hK3rGY
caZ5URgiu4rU9xaxWJdhU/EZuLMcpedw1LL8dUkxCHuqvVcx2KVwt19k9mktL7JPkDWTrqhmORr2
mcqRtvoarcJz9fx7X2IpScv2T7wfxzT31i/SAGa4+1ttxRnms4Waknm0QUk8kY7HMIr0Q5llIRft
3jBoC12+KFFasTBdR5ZtrfGdpVaas67qa3yKQ2MZPGyHLEhGfBcdfSR8BPC1KukJG14yxJhNW7IM
OtW1+jGwJeqERPbb5lZk7GqqMa1Q5d+Exe7dHHh1SQZ+wFt1lj3WdViirW9x1+dQOaXDxSZdV7pQ
mr+8TYCIlkAA1pGme1nFkKY9alZpPTrhgCw2nkk6cUEHR2+FJCwUhDWccr9Jk+N8lElzYajnCYEh
H4hI7eBFzt3L5wO/drdrT1J3T7LzUG0qm+8tQMVuIWxlHWkQ42TwzlkT5B0J+JjEw1wh8q9TvjJ3
mLuMcGaNl/Dhbd/0EyZ8/aYB3xGzOw8yP6ynbkwLe745P0Kana7v3FLSw4QfTjxBxAJlqkqYmCod
bBBX3u5HyZN102oVUm2Od3hagRyBWpV6eS0GDdGf1i+3mp9j6s5PAdUqZvdKrWB6jDmT5xZdnN+J
CV+ucScFWNZStKeDbiUQn5zBMeE+SF/c5BOIYLXsstz0GXQUkGhT+/B2RPg3I9wDWtObsqVdqRuK
vGYxHbnlh77lBXI5CllXT7UQgs8DncfYZK+mNVjM0VbcyNa94z8Uh0UONCd8QlApyFoC8W/5jT3D
rQreMvLmrdH1rppDSCqL0bBXEZVkzepxNlpJBOv/LBaSWobW2bilLutwEUNgqBNyaRP8o1F/72cZ
aOe2l2gEBnxMQjBG8LtfgkLZIZy6hTdId92MTnodhCs9w79vuSYm8TKU12QnTKxE6JXY3TW+VBL3
clwn0r+Av2gX9WapZajbLBQPNcnXjyW8bqa6c7sIrNs0XuPycltu52DmXeLG6cx39iiJxxeAkrlb
WeQ5ddbzq4C4zWUSP3Z4lVD5VJYvOc7qoVxyTOOquw3itiNk453JuSiQOc+csZY7vf6o2Tc8U7Zq
SClwy/orJWZT9+QFAfS0/0HNvMprksGR/Z/cjZZ/yVyoAC0XPsN9VPxrFi2+DdBgpNEb9znILA8/
qKxXnN7Y/6T98LVsHWeEVfu4qPdu+vsTevtZ6rdPn7cjdQmMbLAi6GAw5ist+2pogVcooZyYNPNm
DblYbZrCEDE7EeMKrCxUZPbCNKs5sx+QJCyLoSvupb6RF+otTeAqdo6fI/VBRJt0Wl+Av2uM8kFp
tJ6PItrlOFeoPYvZy1fUkqZInmVWZxdi9XX8rISOxT8DPTqyvIAMVFc2ZlTW/RPj6jlQwh0Mf5I3
jHRQD02KG7OGZcJZefdWskHRRcPb0I5cTY4ZOzNoZhi34LaaWhRMsI6ha1ziAmpH7XF5Bzo0fi5n
Bhl9wWRBAfqOc/c/dklFu5xIor/Hb3lLboHT5j81DY+SbxcxtrggFxWXY52EAD8raU5Ul7rFj7Fg
BHoSfQm7/YO4Z7un0wWRU1hcpQzjIuA2X9R9EMrgeo0COSrRPt5Q8VyyOxogDYnav2b/B5APjA41
3bDip/GkWogM4MF8Wm25OGEXKVmsJahqdgnFb3C6kgWfjLuJKQs1Ib1KWJvAfAdY/8a7OzMdMBum
27chaSmx/3j6SsUQVb6l/1AZ+dKeBIii2Nt6w83Yc64AbROJr25y/Fyc8r+DH2TkT0JpJQaMMJqe
/QmMAs8/cvt4TPOaxQ6tLSrxZyCO7LA1YU48y/xg6K8lEb9tjEH/wrqgSFB06rOba2J2sEJZVFDc
6lefmi4V7tHxb0KeBNUG3u5U1kRYXZ+XZUs4MgzjZ93C7Tlb6w9toYvxqhZa2Ga/x92TQwol6lCS
GIb4bHjOW4G3i3MF76eF8qGQML4UDnTi22OMVPv8oHQZGPROS2k+NNCd0GYum82uhiOsUrB6Cq/d
iIwIQ5FFoSlsLIu9l6ghyfaTvNaDEmeUP488l3lwjcQibNKOB2iq0hMSGVo5KhIGngbaDNDmmQIu
0YjwI3QXrmJahw5H/Sewg1yh//OkGK2cvExdvCtNlXRKb7+H3Em8hdd04FEO+coFH1V7P+WCY9f9
bH5EPKE00Xr6UT8sQUgw1KuQUBPl6xj3obhc8a7ZwKIkNbJNSv2AOp0KpFoH1NtPNi+EmVNOx7ev
z2tBdeq4IZDfwBtPZmRh4kWjMkOKItSQnR59sRre4QjKZnkb2LVxqrtutXbhfmXd2tQ3nYGPmM0y
sH2b+4b1IKBeebINsS/cQ61pDQJbKynfNVCqt2wjfplIr+QbA1du1ThP/8pXDpNMsQ8KHTro/dq4
DON7g6hd/bZAJ3BFp6Wq74D8KTxzKq+1r6Gad+kT0fJiDPTB9nBR4OPVqC5cmfDPqmfksn6TzW3n
+SDss81OZt94SUu1i7kDLXP88sIgqXjTuPyX+pxAbAxSzWwpF5XBfWOAswkHlhvKxSdYgKgYn6zu
AZvqO3iGpsLmrOJhVgN0HTcf6tLijmWvPbT0GEb0VLgyck3MbXcmmhY6TvhoaqHhocRX7fKzFngr
xMfoSkJoN0MH0qKzX8v6gFnHLK8NrrKpoXF5NYK87d1fKBcKbp0BG79PezhnzjM3Nz3zPRE+BS3y
3vJHgvR6hAIjs8rrEKaKS4/3zIiHxWl3TjKaD9U+YJUwmDK5YAv4C4P8TfUDtALHOPvobsAH7q70
2oALCi9fcwEQGCo71a/I8FL/exkDgSbJjb9SePE9ra/tXTj7u4NfMYbsOR1wFJXGrQfk1mEnJ5nf
F8/Hcx+I+Vc/BwQMFxEA5KiEDPlMf+ntFjC/mS8KakteyrCRpaVza9VLKZvaKzbQ+4dDlHbrtAyt
y+h4I2RfpwDDLBJqjidvdYPQ5y99OoA6IF2/2lhiyVEspnwspiYmzc6jKUshj2gmze38BDLJ9vzG
a2YRAN4R3y6Apo5qWg/jtX43ASZbfx77vcLMPr+ez33BlIgjL3A4fkDJlcTL5tNnO32fx+BDxuC9
AC+P2RUXpZJc8xblLy3j4OgsbHE3YMQcdRjHXrRUqN7eIbZw42riQdBbMrKRqhGp1Q35n9Hhd3JV
X4yztWd764rr7Uc7JTM86255YlOnXzn4obKow652gMT6Uf3ihpWbmW/wz9GeHXAQNfukelXWrjtN
FY1temS0RH0lnZtcPvwLfIrufNHTI0uig31iROwKORbmwTkNG2YwFQ+UHtk60fHan237y3ry2UqC
uAEeuePAZWD87mFy2T//6FnLj8nnndzzKY1TK/1MjA6M4QaLUADlj3p437flC1aOSUkl8skMC2Nt
yIaSea5iQahkE8DDmfqDQi59hqCrhmE7ct37WnXtM6wFe8rLaK4M4yEImymC/17qcRcUIMG/sTlH
rF+eO4/0qqBme2mAbTvolA6D6V7cic+nvGK576kL27vv1l8JgiO+9dhIZJ3SxZ9PT9B/WsxbMmPd
Zja6BDYJ4u3C3oR/WvodzUQSDhJZNTJ97RTqx1kE1dSQ4+R6iifqPZ4x+rYwdl8t/YhomGtvHnb+
9N91D8cKc/K4+TqOi6DOQjVabG19YoGeiT3zPqnndEXEQmQj1wYXXokYODrqBJgjsfxbwRtgdUu3
XlhVzp+yCoh9Lza41Db+sO/pVRifHOG0ZSOsm4hizJmIDowL+ljuWdpyVKXUJwWWM2VV2gkMWxNa
o3JC0HsIHdwOl+k1TijGpxXgQg+zx+imt7wODAJHb68w9tY0hz/JurbYojh02ayOkgqCE85SzsV8
zSWOQbr7QwxkmUIC4A8wNFJN3elGEp9Zpy1dW5x0OnpBsoAIfw0/Dclrh2/H9mQaJJFuo9Gd2ng4
6rD3qT+ClPADj2QOFLJIZzfWWVSZdK0UVaBlixGDolEmyA9mfjfOQhCaei8n+sIBjJpUXHyNaj4C
sJL3CgQzP39S1JqywxAkIYgeePwMbscpSsT86D7cUSljw22izWsh+cbqkdYaSylzCu9W1+wsn/6l
2XeUcnpSdH94bmjeGPy595AYWxI54BDlwKhzt33AgfDdgZofTFTfxIkZUy7jqwez8cAiDh/K0zVy
HOS8UK3n1FsVJey7m+1wTNAZM+eaLAKN1fYXIimTuOnvQ4yDccR12PDwLZz6kXrsD6Hre9qU5ICE
JOIu++mLo33gXYgjgfPLrd3zCb6+9xQljyhAZAS0uFwPoGEO9nMr5oy3NgpHJCpFmSA0Qd7aNBCs
TFB8w53hUaOnBxVTJXm3CpNzW0C1824x/ixttkwY/toTxZzfQp2P36xgDiWj8lc+q2ytzJkBY/Tj
3ySMlFOe/WvLUny9xcoRLAo4kiQC+6dt+6f4eiddHFPBOuQsrXuxk1B+udY9Tve/bJblciBYN4lk
qOMJjkqnWXEyRjBBefJLIQ7geCEsSzz1+T2xNPd2xmGW/Jz70xEQBKZdK7rPeoPWkMNjY+ddoMlw
nHczXpv62MnAJ9kbEyPcskKzoJkrriFi60+XoC/WskAKcY2qAUn7FyadJV+8cpOnh9ze3488qELT
lwRZWXSoOiloS679QU4PWYcWL9cEV973CPpS9+TwlbtyPTOgGmOkQ7y7CwSICbknXAFj0gC3Xn4q
dDmGYH1JQiMYQlh4MeAbpLtqoYuCKkZvVa67t5bo43twAB/qVMlKyBYcFgPiF7F3X+YgNujgoCMl
nQ+hWVgzrnXrf/hjRYP9gDHjVBbdDPdN2Fxh1J533ntf4bqlw7o4RNXyFAbPYTaL7qhPLk04KIP3
2irOcU5yVBsS0qhRRwtYELXhBbaq+0d5uMLGCmAclh4a/2dxTf58ESs5Ulgn22uAsCRoH9ZTHBkg
JVgP5vEzZPKV/TMlHZGzzlxdNDGrwkB0gpnOCTyD1Ib7eXNYK0eZ2x2VYDz7vJ+4rFGZloUwwZAO
PnRhRJkrukUTtGHeMN3ZHtS/MC84GNW9xvLILtYym4OABOTC4KV5uYKYo9kHBfUm7PbM+1bxhuYR
LT0WWMwfVr3p/zCNIJAqPSh9bbpZQbopshW1Os2DsVyxWWIbHm6H/10HO2HxRb8+03CL70fORFDV
mgmb3vPwtStuW9lrp9VfjktqNz+tffOl3HylbA9oF0Y3tXMS5tDO/lLXnsI3ubluK0uPLrjjxzJ2
70helZU0Bh6xoleTObgaCSDOTEeyRCORQbej81aaTKtFzwcYxiyfUIwa9PJ/aKcar4ItqR4RJSZc
KWB3pjFLNZU5YKFLUUZMkAIyKF63C1zst8M3ep4yNxHaXYbBo8QBhQsKyv+IL10M4wVmFEl7M8np
HecOSV/4W/TfcK1IRwWZ77PVNVPoPNI/ySlVZfk0qZlABBto3I3OapHux2loTAGnnGKzqTWsU7r2
vjoabwcj5s8LCAb5b4VkxVb38i6R0oMB0lie3fumpROn4jI1JR8SI/5tc+eLlKpo9kR1fOMOoijF
TiW1vbNs6NqL8TTYXsqFbxj4RXYYgRj0RB3Nqu5jk3FVTUeNx75M8p34KOWttoKe48SBGHlyLnoN
2b+k+jNBbFg09dBD7MN1bcQE+69cAidpWao8WRNZUUKyrcQBNIldHGrVj1bZSfwmBBdpJccztP6u
JFJxY9EIXdk/6NcrxB7zzlsNnkrntz0Qj9rHhd/kdCRe6OwDMwH/4e8n6weFpLnl7mZbBrgauDJv
5eIXGVFUTSdybtUasoq2mHAwzCotTY8CwuuYWmPFeKTGhJh3zzAOSe1BKY+8Ip5Ovu3ZPpjTko/a
BkW0zck6z4vB2QkgfnaDYUxYS9twTpCKTwkSpIuSWFbdAv/r+hRk8ZBDa7Fevxzuh/SRmtVoi0K+
ju+0Tm6/tWm6H94RxSDlZH7UaxN12W+JFd6nqfyqTYyVXB9e8N/ydhlPk0mtJpb7FO+ECBP9IGBN
bYgAQhg2JkXHBX9BJmj0vlFa67W0CA3mQGLQ+tyIDsoi+LLzpG3tidT6PMpPqQUREVgAurBC1npA
zXPBHsc2dDlWmlf4h3zhRIw+xNwkjxSbILoYBHhNntn0dLF5jOM0/LTYNs9gKKzgte5MUx8iUKIz
29nqila4PsECPimUW8XMnjZt2RdHk+49Qn3YtbL52xGh9qQ3E2C27KtTjTP/KPA+9YbNNXZrqw6R
5g59VkMyf5/dJqcsL4PrYbK9Y20HvN0BqLekKWAx7zdbgmb/1dkMdaiElJilbo5OC5JWJ5gzrbb9
pmjSrwgV95Cm+wApL/FTM03/fntRsB78nJmu8ev/JKuS362Ib15lO8tW2BndOEnVRmf/errrXQYe
V8w1m+Vw6/1YG0B+IgaPyEsrRz820d3F0AjvsqGDdcEPKkkXcOT3zl8hLSopbETpuke0/dP8ATs4
0igBV+5SixGJmDByIrahgoRjjYLf6/qZASAxvf7dBcyqH0ze96Ynw3V6RFgyxIGBNXlZ5vZ8uHYE
CsLO9MqDaz3uHdCuz1bSRai2V++UT8eqwfxiWhCYAc7gRqFLmMQV7CSzicTvXfO4Fk7uYAiJhH0u
YT1R+swsblRTBbDRVo4KpjJMJd1yTjhrshrolJgH/taMeO4m1fl5caxf9MgbDXzZUcwRAj3d6iF2
RQERYP8Rik6TJfUTSB1Xr+XYVZNlCuiP6zfg1a9yCxzzpEAakWgrFsZuskxB863Sz315JxPiSkc7
MPYXwdO+m15ODRiglMklHxALiUF5zCsWeAywrpnVgbBmqddiz2513TIO9NHP1kHIV9smqGfr/zfr
SldoGm9U8glAX9vLxIiF7nDzbGPg58dcK/SiWGVl7ezeYPXpaydkTrAaOSFx/kQAmT+HTKJ+bzU7
YOSXxq3Geh+Vu6EgGzhYh6DboQCuuSXi1A7ou7aTm+l5bjJ+Z1O7O4vyx3mgKQl4djyVmHtmEM0z
eVj/OhjI7gffkTm/sH7NPvguCsX46e+pUO83Mkay84rFOOWFHCtNmIMN4WV9MDzPbsstwgdl5XBN
ww+T/kJTbkEz+KoX3h+TP+oUECcwAh8nv3FCjRgcHaEDdRsmLEnHdzbe3uGANsu6HXAPoUBp9KJR
VyZ2zLev7jCap2Ttq+Kupu5uSfYhC65s78j9FB8ncuxGqsqh+omB/YHw8zt2ZvGC69qxbdYv2NjA
LiT2x1vGOQ0FJ3EawO/oET+JqiBvsTOl9OPjzNbMAlyN19r9lvYPYGzLJGgyHT8FB42SwAY8pbT1
CLo/nbx7L6b4yM25zgJvIazVN2FAzp7Y2F7bI3OmkJaHHENLoqz9yQYAB27VdwMVVOGCcBLHRQqx
SL7xmUa6piOplbyzRIv9kedo25P2QyzdWbyZUWWKSbcN5O6YykGsO3jB0YvJtfv1bjfneRA4fWe4
8EW4u3jRF8MENE0GvW4MEBYjBiTGm9NErGN5MIJMH4zm1IOVT9PJCr/I6KuKRR/G8Pp5tBqBNNg0
qlkryeCe7EkEQ5CeXMgTSanheipJdA6KWXyjCwrcfk7UOWKoyPeHaU9fwyMcGXRvTLtG2tER62u3
0tMiXXHwXYCPDVQ7pUCEQVGtIfOoBSmbE8oJCku02CspcTuWfEPPs9jXyDkUq8b68zG3l4FN/bEb
dpmiIOQlyx/RMFVIhakGSQZtbUXXy9ZIclxxuSEfraa8fpyda1zmUOVYFhW6ODRXFk9IfN9S5gI4
CDHe8MA4yOi989x8unpOirYaGElTJhG9lISRsCIWr7ivZjDEGOoGbLrxIE3URxj5estHT6JF6Obw
kLOH4XTYYtUty/lUCpKUC1pg96vjzEGjOnnN5fHmWlx/5Li4IWXQoGNFHUothb5MLEFk70YapUmB
o7jYe6EBfL53Q2Ay0kXtlz7DxK6ro2RY3XgJOGOAxwxwkp2SAjraVDktBtXgIg+HK93NPY3nP9aX
mfJMqYxwKtRdxx04RKtk+qmjK5Vwv0O0D2/AOEITRDqqqGv6gp9W2jizSNwVI3/qF8Nrdqld9WPQ
AblsqOD6ZIhiiVo9lFb2sGkCQmQ5tSamfgCp/tEmAYNMe2RyAjRrxfcEo5oHpikQ1RGOSM2eID8m
NEqUdVRYO0DOL7wC6ckX/pBpImOk2ndEBLpg5wywVmRZIWypT1DoV8Hwsu7Ek2n8Hw7bF2ouGxj2
c8dbwe/2UFKZGUHkepa7dEoU1a6XqHRuvR9SJvKk1gab2sPkZZtTLyBJAS1pOKomTpf8o05PkllN
vl65KbrCshvU2YHuXI4khW/Hp9J3X5006PmiV45KDk4VPiznU00ijpKoPn2JHTQmgfx/iWbVdDKl
VaSdJ4/WMv/EMDMDgutT0QAP9GsKrNw1JL0xU6vS0dUc7J/Tr8aE6A9w0uhC7JM0zrTTSJKAhxju
QnD9mLWS8ZdBjdkRbL7TgiZ/z2bj91Sby7Dec8trz1wt6Tsa5OJ1nMS3U10wRn4Z3R9TZwEQUG/D
dK5+9nP0ESb241WjKpe3aTdHwYzoG6gHqre5gH9qcDWnA1fUXLEhoJQCUtF97HSP1li8CpKVks9P
EDGYUgrNWi/4SoGtKPhlsy6U2cxd5/LVzts5rUhRPQqbUSKW4ZsdZ545esd7eXM21bkStslH3naM
vabC3Y7pttYo0+7UMaUcB5AB0+2cHHvURTNvzPELmGNWFDMZTZiJh4ts0sjyMx1Pm9d+mUP0Gd+0
BC4ULElaznLYhLd5o+SeCqsxOC15fY3qjEiujwm+w0r8Q+b3bkqigARDzPGRO/I/5zqQyKxURG5y
9SUot28spk6uYAOY4dJkXuL3R71XALV3M4SSQxTkzLILfBPafVSZgZsK8ou/kHCyw5XJsJUEciW2
gA/LDQzWr1HnQCLZ+5DMoP/ls+en7SCr061HvCnLe95wPkk3eayUp/KiR8FkMv47bAuMocLh3t0u
IG2zd47YuP2oN9+hoZBcnHvjLmN5ps4bgN8sEmmtk07hFUjBrlSUpEGY+plvuDUfaKyL/99DoGQD
2So+F1W04HEv+7FXfL4mJbTxaoFsfe7462vEnEQq5WRQi0aK+Z2TJVMWceZjmRpxZSc5C4FugmXC
br7QjaPRxonBFflli0f/qBm9WKguCcB7MZFO/OrxIErzVB5tNaAdXAjKmEp58vEQMdXn+/LMO9n5
H/cs1nbNKOJ5jLFAHQ7DPL7STv6rcell7gInEB47pcEya9kce3vvWndgi0uCNbeouNI0fOTHpEZ1
v8Xe/M7UFPo+HXXVn9dlNboxjxXqr1BuFXFzoNgAa0xaH6eSSBxj0wHg8rfSWynfLIZyfT1JnaA8
3Ya3CgwWoiOz/PioMovVAqPUyD2EDe/Box7foli9esvwrXoXnLWy3u+HBfFslbQ+wg3r5tZEiqMw
4ZtjXmz3ICdpKqlmfXdkGLbdjZ9nOfMhuWxIF5fWyZhvcv9vYh18lgMIiAUGAOYGc+hla9QOn4r5
gLQW1X8KaGsNxgPPK7siX8kuKWti+9AdAYUilHvcUqGzCGkx0iuoAw6RmAagBgcebrfLw3SchOCq
bot/h7YAMjy1r0o/ovR5onODK5oygc0LDHZBWz+nDiLVEhw55DWR3+4uXKk/Pa6sPbOkwKufio7U
rfGXpKsIGL0zqcBf8SCKLdz1pi/rzp6P07RRAkm3bkcRYZt4/YIN7CzN9qw/g7nhzq05OeBdIe+E
iFrD4rvLKFoDkQ2o0bK1OoV/7rNsAtQvcow0J75hJAxKhDKjLK6Wt7PM43LSa8ZTqEhwrl5/8x0a
zh0W2UQn+2DgKZ51FbxXU42gg2+QBZUlgDHXdMwHUp+r8vybBtkh0zjBS/QKUQkgGFtsRPj+ZBlI
vsaX3vRZBOjqYy2l2fVNyya78FR9O/HiELqvdbGQ5Rncx9FPppgdNjdbb87B2U7kj5xMKihD7EoH
cPx/3SjtgILI6MY4lK0kFwoETWMe9ZORFb1rQvha4kUfgtrwnqENCEwIxddVLRSC4/+HWn1S+AIq
vZrYwjY1rX0aGz4KZ+/T+XKTyS6QEybaxzORQh91kXKYPPG9VZlaF7EuqYeLRhlupjmJOS4uaT72
E8YRzcncSFHaADGAAQmSjci7t8+kP0NJ8gFzYOBMgsZ2f5OBCdDvAPiPT6ObAuFfpqkl0LUHE9bf
YEJmy6Y8QByrddCsQY6pWuoqQKj2EnHWJ7f5MZDS34sqIqMg2IMB+GH7Mi9O0eTcucIi+bq1WWZw
igImcbA7/Hu3RmA1bRep5LCXUEyMywFJldaqqmrM/zqKCdO12xbaSSypn/qT4nee4a11UM+3j7Nv
N6PzvyINIzVI8LUSxIVEGOnpNJRvIZ0nxIbKCKzFTTetw4krHKEitEDsojnu1CEwFRMN+xNw8OyS
HbzmeSrE68gx8Jo56DJ724D7Z/MmxCF6Nvzw5EdSVUoVsLIyir7d3Axoj5OsJZ6TkRNG6wgD0FR0
lGHaQArSg8a37L6CWMjWoVR0iayQhJUN3LYAZphT2IQN2RTt/9u1guB8ExvGFTc+x3Yb5vm6AG0Z
S9BABhrWBjF2MOgejh1RVlGu9geSOjlbi2/vgzhC8c2uFNj1dcODJpdaHJpVl/ZxtLMJND45sn5H
CxI4xbfmWON+0DbOPB8WVz6f/FK7yNq/+lS3JmB7xEtHQYejWYuukbWiSG9oPa9KSfsKYfASQtj+
GrALc+o+dRLcfgnxOPvfYinnmsrZ7wPg1iXZmpBpTeLdd2VeA+S99SMM7cS7FB8f5Jeei9GuQdr0
+qS++Q8iqN88bMt8xEFy7vyvLLbymqfGQZCoSMvARUdLNNXBvgfOyyCD09+CNJso8uMw8cgiaZsW
cGzFjvCkhLjC33WZMRKSKvM+8Zg/rX2Ilh7hc23s7aYzUI0O6PwUI5MhgEeOO921FS6aLMlUlvfW
1lFsDYpQYCh0TKfmkFyLrXiduEwcCJqvM+V4uJ2ao2om6+iRBarFdV8L7qO8n05OTaIgK+hAlUFV
ix43HIN/m9KRkItOmYkbga639ETt0wuXKjyORli5/ucEtacN9lgXzI7yxG6QY3Ol64hgbcUzr4oc
r1WOTiuufeRMhmAUB+XbDlzE+oQnUDgPmwfUonX+2tdi+9BzBLUmVy7eGj4gQYYEN6xZ/GMRsK1k
oTfjABkO0MLIiYVkbqOaNAbNkBzRzHAKNzZeL+GbfDaCa+YFKrXRwtxYzQS3pj3RPa/fBgzKFIIP
CNOSC7VAhPZLq8QLB+vv+zz/MuEeFeI/NOEnoCGquMGHSI2K0J9TosDyIOuXEEF2hEsWMHusuJZp
ojAoWn72Ovblx8uTNuDuhHyrtYZ2vygArlZ0UeiObURe+W69Jm9+cDVg2jRppoXatM2s2FZac717
i5AZwenciWNrcXqwY7fGh/SjdPDudpFG+xWueAv4AWvY21S95SfUG7XEiI/dmgF+ZZfeMweFmlZI
sya1kbNogViyANgujCzyIhQHKL9aIhtqOuOZEwVLSGVtFx4wIw1mCpiy5GVZ2q0OzOmMio1kHjRp
oMHEvXs+3kpFl2R9F6ZXVHCyJqNTL7i1M3AJVP/m15ILo6nnFEdY+MxjkeA2T/0gtlRiTLOEILoS
t8ZJDEY7yu2hBtqfvEpBGC1NkhyvNuqJYEmjWQmoQGG6jF5aAYRm+TKUJj6n2ksrfjQaLYFZyMHk
XEMwb/6hZZdH2chGWgTo4hynJEIBobZXVLEctWotN1sU2JtcKME4NT2/OzsuLo7869Ys6JZCOny4
CZKsrCKJYTvGZlEujM0UNVbgpQjcKIVBWg3UKQaNPZjHZVM07QpjZJxj1OSXdzHE3z67MiP9JEdM
POMHJHrnsh87AhZnCiY/jIh/6abKjsz+DZxAu10sGs8j1OyzVgDndEEHxofayML2u12ADue2dIKz
APBJLr0zMAQ4TszVP8OBQjtqELJcYTrlOCLgpWNKBPwzkbtmC7hqSXsdNWgGd18cLS3dLTWchksT
ayFxgxcR0kDhsuiSgap6Fs3BlQRaZfXzDJw1Uxiv/L5tCK03BQT5+Bw/y8ITlfvUeRFkPzOtSf8C
wUh4bnN53ph/EVbwRL7Yuk3NyqhqFawxQd5fZBYCT6hcbg0wYiFGJe380rIlIwIcdT9ZxT7r7c+g
sRnf+JTZ+t1Hh47xcXDbyVNTt8T7YKplcM6qrJl12aeRbwmj6HnLDm+H8RjiDeI4wM9tLPV1iwNa
8hJQW6qLAOXC5tGHPsj8Gfc9MJaj7CFjgYL6F8yOMCZ5XAwLhUT9PfptfZD4ETY4vy/luM8pQ1yn
rWeLZVH9YMvyb7NCDMyPUl+OdUemZKG4lSnWHd8FC+SknbgOX3LmiY5YhOPu+oAJr43R/XBjiEV7
29o04+6nlPphTwFyCAzTFjfS4LSP6c+rdwCofNeOtmToRSduYJvojYfUcd9nY/Ss9Sa0XBBO3v5A
7flvvC2LLZmwqJIAuFz/X0k5tedMsiNUGfbWs76EMLu1I8w2bLiHlZyvYe2zGW0MD+8CyHpXLLM5
vPnBZt8kEXgHWBVu23nXJ3xsECtunG3/Tvh4j4Iye5Cg/2axyb0MMrZZHX5SN+qZkEDnTw4dRGlY
p7dyqRjs8iKDTUy35gGgeI2THtaRmBEvALLYoK7mQops2mP4Guq1i/fRNwj00P8v1ksCRUJeHDLh
6yn0mj9Y1n2yVxeW3C0GF/nP+Z05tPqjPjHmU5/wzjpVVNCk1ddsskZjXV3FpI8h2A53ajgdS7EZ
ZY8EM9vyZ3SHrhkh5/mnGO0wP5KyqsiUurdQmDG6FDC7GvRe5n93ycScNvBbR+AYxanP1M2lrpkj
UlPXD15uQeqKU64y/B51fJJrs6qhnGIAxJ6QYEVywWZI+w3Tm6nVOn0k3H1WJ5a/tGikOqXuYuoE
uotnte66F4WJodhE+7rs9AL4Bp+rdLk54koBETlFZwPQrXRXyxsKJb4cKOEiVT1M9KplmjRpZpQb
F3wPlxggcvTmttTywlpeivcIfjoS8LdN6k/qhmeEd6zO3VurIgr+g+RMcL5YgJYJUBxHpCbhlUh+
FSKsvQfd9+xxHJ7vmwNJFANpECb27NRASnB0DqMaZxL7gFpivvr23pjpxRVdxIWAhUsjHo3KdQE+
Cz+TML21q8pXJeubbjyPKcvxsxJF9oGNHr6dvF32qMfOxpQ/gZESukg25zLs7sAf+krTAaeMbsYd
aP9CgCEUxejwkPPiTL5gTp+kPdBRB5S6Uhe8vJi3q5Z9Ozojnwp76v563S5NgbpCNvrn9duLoBd8
VvGOEXfFvVA2iPLGuAIQc1OpYSWFXg8uA84OuDvRDxOZySUGykoc+nROTMUevEkp9NmM6vXCEmRA
yDA/ZvEixhf++q7hFbZsXKxaAr4/YXuNpaoAeSToeaEtKjE/DMr9nrNnjBzf0eY6x35Gozv1JR6R
uGamV5mP9YSMmzWFuPRUr6UW9DbJnKi8byzO/wrzppwa0gT/2M/pYkwNgUzscgLYlmo8QkB4StjA
bhnj/AOIzxRXPuQHt3eKvoJxRPOdLsI+htEbR9r7re/40ZK0o9cnsYKsNnFoyCg9hej3ZXR5vQ1e
r4W5WGkiTooEHGMU+r/yQRcadL77VZxVFpilJBcb8Xhweefcvh+vtHjxyJ/AR2NM4w9++FzrbFLr
KP+ZJkabdB5c9mZpl+XGGW1l1ypsUvxjqRomgOZhH0lyl70uY9sPqdv1HSSLTz9O2SOkFx6GX4GZ
SiDCacwIsRR8My4wcdErrZgX4PWn3M4XNavotUfhQVLyhytRaXBfXlbGoHNm/0uMInjZB3+jCIQ8
WQWPS1MRDkqHHD39BpoWJya0y6g8uP7wnFC3Ohyrr/UZ/CKWnF3TA8PPYvzetK588Kx8lU3Y9teF
8oKvlHAqvYSHnPSxBX2+agjqc3cZTLWDwnuQffNyszNK2v5b4W5jGeoH2GQrjzhGrCnusv0haIJB
1vISP23s+vS1G9wMZIisGKGiUZlZUuk2Hg0Scao6FjOOVkFlQd9A7/dh/tKGFcJIp7AFe+QdQOfH
2rw0Ablhk6/L2Ez0IWKLdg4/mJGfxgXCKrTfhsLhcHNCt5n8fKFkt1Y+S2IZnM2Z4AQzqHiyCIxD
P5YABdjeMSS1PZeAtV/VCdHhSAtd/sKi/0PcY0jndY9HPAS0OOAl7G9yfpHVzNuBSAeTu2/3efIJ
lfhLTpi8SuxVMUd2s2aGgLfsoRvNoCcUxNoxG1Cawnpy2tTaH7Mk4QOOCRh9kPJ/jEOjD85qJ8cZ
y6+hdG97W25QjtoZ+O9/++Ba8DWK8pIpgEB4NuDiQG4vhgilevlK8/4rKktLo4736zwcJFYJTMfB
CWp71I8NuO37oG1A5QUMLgnkjfoYGNjgAJ2AbbJu2ta/1J34mgM82dkjWH5GjnVUL1bzPazESIS+
HMLsbIFf1pet4ttcPh+bU2sIw1TDq/PJbPxwo11BMf5HJOO/3ImWhznPg1knzvSnWzCuOHCVy+WJ
feCgJnk2jddm2AYezzkjMHRTujAWiQ/EHdPuJz793AbkK8y0dF70aYoGJkZ9AJwZgIsAmYP57X4G
/tecvixhek4f1kFV8vvsgjNeeMaHsJRMyk83yMFazMDlB8gdcQrKEvw/62q66pJ9YqN3FCCP6qX/
SnlRRDXR5LN3S56IbTEpdQK7jWE6hE6nYRlaKZkZ5Sgl3OqaOd3F/74vaOkG3RbmUq2S5Udo0Rfb
Yj/8rsQ8JnKXIbEHadq/1jZsaJYiWoXG3dRJsBWshFuosHrn4TUDLmQjg+z6LMb2QpHqASKeX2aY
kEHYCsVo76Vx0wKxkA8CiEPYevzt5JmIXVm7/8IUUAOdTZ69QGEJFky7i9iTFNiG8HOa5AHH8ysf
6nCP2DlsMN2qSroTa50iYx8GYAs1qVUQU35RZ5VD/uwEP7HfzeDkgI5xAUYolxK/IqQLLbsD2PTq
xIJprRUHlIYF05BhN/wBbrSldV3Zjcy2iLGRyw96h3d5e180194vTnuSSqlQWgE2oxIow3oJHgmO
l1XTNq48LUvTOphC9yIGq9Um4pE+8NaMlSzoYItayF7qbc0Y311CqMyJ3jJZj20SMnyKmGBjm8nI
3ta4nJR8WquLXgj08+SoBGlZHRkzMR2EWkjv1YgXIHBWDeQx0sMNi6Hql0vAx6uPU20jMnV5lmKc
F6SuAVteg4q/4F7sgiEnEqeln9nldFNF3+noqwRYAkbOJCy/mtOXDk6xEOqPmaz8S/i05EQrKW2d
JwtYcNopCPI/0N24uRqTz0zJKClqG5cBBU5MUR4bS197Sl/Trfv2SWm1XAwHgIC3weJu43pZmR8P
nbf8SZwltzCQtt+xVIGNIlcvVn5xAsdYOVObLbVjsvHcq/C9WvYbA7xGsyfmpIysMp/aG/zq+3ld
upzqbQcPixh0dVs12gA3VqY+NIWsJF2CknhQ1dBeRvzt+mRcd6MZQEZAcs9jE5IkldGb6oMV2lJ0
QplGqN6wIkzk8UnQTaDQUJY3/edTypO5j8v2Zby7oAqu2tHunRcfnSsiqtlXmhRl3a3oTMGlGHwB
d05tQNkUg3AwdBylDYKDAGN6tQps1q85sVaW1daEBaH598nm/9LcRCBptTKJPIbIOP9AJj0haEBz
rZCDDehHOoqPHUx6KCnJf6xNuQ/OWQJjgvoEIUZnQ5MZBLVpOggr+h2ltTm7raxEitUr3lFMlXRB
PLXHWyAA8HvASlTONLKbzzyr+tqgZasbQzcsfHmL4Cmh0+yo1AQb9qQVyPQDa3j8y47ziyT2PCNV
OcnD9oWDJDS4lS0dSBIy857P4jOuwc07PzTBzVzR5CE8Np6zCwvl05aM8i1KEK2sWf5f92Hu5MXM
8X2Jx1OYnDnh/Bylx3vwnIzSnf3Sk6s/bgXt1hUXmPAuEZzVSQ7PV7oV87ZMRMOUSiWmHKUUjU0y
e0cTBlJ+yQKc4GuYLSzwZcfJLAdUp7ydJMki4MRSfdn0biZXfJIl8qtI3zbJIQKmfw418xuo2hEz
eY/Iw2o7cAlKEAZ3H2fcu85LWEDjKnkP1GGof+gUI7ttaHGte4mrPTcNcw4zTFId6yCuqc0FR5Pb
kRfevjAY/kGONbi+rWpPVXP867dx3m4mANj5PpCVS73CDYPFo/HAzLojigVxjmUpWVT5lRcQ9Axf
qHbVi4Os65wVBipgnMKuWuXexHbB3GmZycG5hxMh5W9PbThoa0lBQce1Z7SHiurPx84/aQ/yaol1
28L4aYEY1ty0OaTinRD37YFGUOO8rMoZ03UMGvHZcHWXC+dYEmromXTeirEQyPgzJGcH9wQIjqo6
Hvn45nrqXiT900RxWcA6ZVEQ5exOMWuoBv3/sqV7I+6JqrVqfxNrQItZdIma+nzsutBkVpa48B0S
mHfdL7I+rChtQD0btS5UUTlWcPSQZaEVDmWJZn5XJdnz3JyXmaesV5UMsTV7+LOtPR3S/2+Gv6VM
S8SHmt6mzL3Oo6s3XEwHp7Hvslbikpk/35PHfzFy0+2fu478ssAuoEzCYDvHNKdRtU1TTyqU4AYq
x6EcntVDsvddeXZWQyqCFz9fC/iLNkO1ImuROwcqgK88HZDPUjeS8dyEVf9zztdXMufR7MXdNq3W
pwcsPXSZKHkRRtx0IXYqD3D3BBAfmnv1eAtXwsUt5vPJ4rpWeCNCXNL8LXLg0YO9Kcjl93sX5Pnk
wgsKYZYxVZjFnAoPQzefFcsArbo3yr70yOfHDVCsCMX68kW2V1eLZx9bjEwon1Eoq75w8y3KwXgl
gfFQ6weK7LWbqRBv0NxBczq1/PHdApnb4/i4rdfJoebxR81V5xkttjzOtu9+WYBPxps/U92M4ZBR
TFHFxMS8Td+AXQxXSO1fpyIj4qeOB+oHOxe5jL4QW6ePZeaNVy4x+MGoSqECybBX9bQ/iNGh6NoG
2xukXtId/TPkevTv933VadvV2bHP1OD7pQZBahYqONtb0r9dGZ26MnNFFdc6TjIvmYNraT2NcZel
XG/Q58kFYeaUgPsxdM6HzSCdf+U4pd0OcgTBxUHXy0gozrWzDh1CVQSYTXVi3bmGXTWhgZL2vRlx
aIcgDAQTr92ytpJNz+SezAynpfHrdcha7MZhANE87CQxIPRoR8DLTIl21c6spMuKGvfJvZejnjyJ
vf9dhjEQBy89tStTq3zUNj3uZZrMdaHASVwUR5Qjpw+ydsTSa6ReyPe1NYhvwyxnFPiQoZxNlVoE
AtPkH8MIvuuhJmsHcThBmP2MIV86sCdloGM2DK+VN1CjKyhR5Z0z1iMcJtE7VNfsjtEH7PZaYhhx
Kvixjk81nK346KZy8qhQU46wjfh+GpbYSSffqeDC1J6QzUNES4dumBIlepnaGxFpF2+4ntlH+o91
wjvdXoNZ4BEOUQIFur0L4DDi/MrNezMxL28qTNCNRbr9fOlqkdbs4RzhIXapOC5oykmNkGZ3k/zX
d06NS3frUccP3RoFhN06QzaL3i5ru9d9hH/GxCU6Mt0O5YV79SFyNJv1Fk1/gdicArPwAAkMaOci
G+OzjYeind1dp5SpxAB4FrqoRFBRt/WarNIUwmuyA9oUjdO2NgiBKaCoaE+VuCpngZF+RA3ro+D0
LukOpibh09zshIcHwl/GJURgE1tuuklxrs/Yg9jvIlF13zR3jod8lJttrFTRRE9wl880h6Avz4NH
7Sd20+QZ/mZp24Z1lsk9IloBHwzVioZ1u6yptBk6kBNHOY7XwcRxydKiZ8wbSS87469mO9djsQ1h
FYCRtmwjgvxAk2iCq5QJJhvTuD8KxaVSHF2Hdlh/d159jE1op0LERRa1fgW+glEJsqnpWz58cfZa
XJDnlJOHkAa3JnPUfm7awHfLQK7wTnNFLhJ5iF1r57Kt0F3D3C2WC4j+IKcFlwQcwawPG7bF42Lj
yebz40Z/0fy9nEiLoJ40CcCe6vG3qMxsVVhcwmK48KqrkTr6auY/sr01TsP8tzlOmZ/kFHpyxNIY
d4+8OilmsXz1Ar0XLfhiTLREJqhNhL465rYfvwom1JFyejcdhQDABtQAbVlf+ggPM7+blNgeayzN
oqIG1NmYP215GtR6gDQ/se8yUBCL3xREdMX8pAv+AXEG+GgA/4YT0OJaTy4kaQVSzNBwJrUVYzVg
n+jN6K26AN/v8XUPB0L1zRxhyGgf8KBGgBtGFqqpMDTsdfAPqbfkUtwe238C4ZiRONitaXukd3u3
IuK6UU8stNpqsYdMgsmuEPUxQsrKffhw1mgR7OULyP5NVbDSLolXRIDqHrOblU9MvhUIjk2L436c
mrzOIaa/dT8NLQ3k1QYwbhmc4QZhyQpSP9cps+eOLvLkuHaXNx71PgfidT5S5tg0fR2vqpfP9JV3
md2NoTnPn87pSrZgtkJOur8vUUsVsmdoGhiOzKud0FmvUeXqHV/uCQ4yK9TJuay7csXeb8fB2kAB
P24WtwGO7yuxzJpF9ntrpQFQZCe9fmtUtRFTmzzC7YJVpRUshI4AZ+cn2ocfRB6oPsxSUAsqQUTp
LFp8h5OWz3tlATfswcXE2G+CmFTkw50f3kH+QA4VoQB/6lpAPYi85aXOp2bRIJ+oHjtN+5B4dhpi
x7KNJi502rO7DLWzbFGOgBRpdvcRdcNWuAinONmQYVaXCPZnlaL1jA8d7ehgpSw6OVJfSoYuuIoY
VSXjRlNa1BGH3bU/LQbrmorrMa8KVGtw1T58K6+2mEf4+Oqm5nJUkrZwCO5cS+nCoQCvYyGF2EGv
iL/y3hbdtko7iiuMQ6OJmakzbVj7Ic2iJWlAN9Me7364XuPSHXm0gmGbtkmAHZlpPtClNTF6MpsI
0yJLVWHXIQk0K6xOI6R3UowzBQlok2XqlmV/A+h6Kt0PxQWj/R1US71Sut9CLV4R4DepsoPY7b0B
kiaMJFmfa1eHivhi9IBL94fc1s+p5G8RKPx3C3aS9D2A5croS8D9ZM3A90ik9lWFioNzxE3ZTtZa
qxP5+JWbC7BGzPeinhGFbknou/nuVnsyiEarJG7L2D23SbwK1+r2Vec7M6qkkpb5PuEaHx6B1IQT
A8uJu9IF8PWXhuritSR6wOZrGwdYrJ8+DwbYpZNy2mzLT48hGHe76FG9Nikv0EISrU1A5i/YdUdj
XKfPfg+hzWeulZyjXfPpHzPoh3yxzHz+cFRbl0DxMiRyMTp+XvrtBIJshZch5E26iLoov891y/Ux
z9IgininPHW7RHYg2WQnLcZwhz8cSO1WvZxu9yU7VoiiVa7Q1pR0Z8b+w0ON/5xyo83G7fQrj3tC
TG2D7EIWQ/FKs9BXl7oiWv+0EBzkTrYKsXZh4WSd+6DCPLnVrp4qzcBmzXFekNeiaHxyzfn5AfYv
rc3kD51gunOfxlzNgpDn3bXxzKiExcYVn5BGTtdxZ3kyXZKl0+vplE1HYhYjMDF2WI/D8D1NTt7T
B8+pr1+kVX/V7IRQe9G8+SVQ+7xb4thViehsE3G6z/wVCnGIA2aQAKKZyfcGhRQkbuaaB7qx0KZP
LRIXcZ0nPRqryEO5ehB71D4ZkiNbZm5YIkMXeafltnD88R7kHHxL8bgiU/0KgNlldWc83XhIkdZM
by3qeYE8YZWdEgSHyVIJ4WqcmDXp1nS+gxtM24e0OX7YoRAqvseuUHVtJKzKg/9uTrjy7ttUfc3v
lLf7OfPKAwWu/ZoVaaCyM/rlWdYoNygjAKt4ydseGYncKf2R1SaR8/nFe8ZhY1TW3kAf3Zv5q+RD
4GgjBajLorRKxN07R8InoDLNY030rsYQX+sAbDiD3V4kUaVHwHiBA+Ay3Mw1mBvPwoAm6/Vr+iM7
+2YgBFMpLSReVMawNSVk1CzMlpXNQHsoLH2mU0MqVgJqgLjhUc7zRveXnF+EIr981O3pCjCN8gRs
OiqYy/7NX2JeqJdzVzTu4RTQwxNsDhLDJsRyzXhsq7dhxCUqRe7tS79nAt/YtY23/5yppWwoKjTz
CI6STU3iu+vCKEauw3JWaWLTRyrgmJKqJQtjeI1SroMyUFGOPbEBeqE91pci5wIGis/g4p6AQqJ7
NsQ4QeCIwlhJDzUD6zkVp1wo0qOtgxSxSEhjiF9ep+wcnKIJ3NAnIZ+zVgSa5ls8DBx3jARsGJYn
+JWFPkj/x9GZeso/Sb4h7HHwzZJsIO46+k2B0P68VW+JHqQeiTUqOlb2nQkVX743YuXdGxvXMs9r
6gOhOVZMLSPu+c/JC9tjLLzez+3rf3ZXm3zeumm40I2geWEXBK2FydGCw2jHgoBGpMZrLehWSWD+
HL0ql+LX4kxBhrc2l+IgexW9ZCax9zmaCqgB2FmrBaG2jGtZ3nxjzq2M3FDw7gvObopZ77SXuqPW
aMdVB9fKmBL8k6VIWwS64GgT2NeJIh+gzUZCSFIsxHO8hSNjMfcJ0sKRXR/pdoj/RKZEHmCACCl/
6UiyKvWIBn02f8atL3dScdrGUaX8plHayHcxCfZTeJdlQWQS2fsZwxtEPf4lc1V3ENdzmdSBcgxZ
XFEOpFVw1MXHPXTe85KLMcJrQkaFLvirIe5Gel2wYt4D1ATA0JToMv84aKpwLG9XzXEMfaUCQFdb
tymGKBozNxDEoLtflj84ExCsFb36sVjK1IRVJ7Z1+Scu99eQ4K/dvOISt9SFpyvl2GOW9v271XSW
oB+NwbRuD3ub//8AGHpJqk5oVYTIR7Ypnp0OP5t63XtFNQWZ4Vx2ZKQOGpQcsCYxPk67qMPVjOru
HC3jd6rFgeCQ/GsC9Aerbuvl+ksQrsVgY9Fgaf3sWdFipvBMKvCP2tqZGvU7qTRfuniQgNYA0SGw
KIVxhBsZreklirKfI6Mo4rEMiHi7PuKOpc+GpETAEpfVFb3NiBAlkFKHUg/S8oAjldTdDmd2H1xx
vDIwKC8lcVsmDo48tBpKB4/sSLyNLd+22ToTRJWgI/zZy/yKKyZR6YmEctP2gVGNoaX6NQ0Mbo9X
k4DajuxxU6Qm0dx5PjFK0ELzbExe8pMITdpkThu4i1zTI0vEu5yWFtVIfO/5ZXc72+hl1Ew9IlDn
++7fhsPXfLE+dwvOUZJCZelbHnePd+Fme/eoBupMMWIJWZ9s7dLer35dLVgLy3lEJ2AZhSQxNM1n
HxmtO/OaWJ6wOyE7/ClW6ALZ5OTsiFweiWUvW5XndAHWDOhjVKiuqEUkFc8bnzpgPv1hcrVuVc2H
ddz7g2RCyQFsXOv99uMgMUJ1bDbHGzVkDD+vDM97I5Ht+QKZcdzHkufHpjVyAw3VvrZtytUsMFYI
9h4rCFlpDVVkkqTbDri0/OoK+9D+C7oMdjv77JsQsccvZTVFzD8117FpBqA6sC49sUqoU8hbDglb
hjQp0A8Pa31Yt6NozQZUMX4JWJUOiJbrxIcmmzDiV2v26B53K0iUzxSqm/lZmtXKKZUGxJYU68HN
pt9q7VyT10IdWwJ4p+ee+LHbqUaogHNPvJtzPAF6Nu7OTvNduoeX5BCIBl6wtDy9C1L+LHuv9+Yn
pkHil9VlXLoiGOurIaSPvIVgoHsVzjb+yp7q3hjG8q9qkiAFYnJaj311iMYxliLf/q3aDyjG+BGU
QT/jP6tzgH3GcB8xjRYB2CUH+okRaCVpPuRy2Z36Gf+2ylxQuAFx9rRW43gt4+c8r2vSShk6jhda
W64Jh3XYzGnWDLgSX9vbuyP7Mraq5aGTeKUdZIftRVHoq6ikd1U5nva3+2TsUNLJHNs4+L9vJCBu
bGqpul9Mtx3H/QX3AlCiikOY2bqgNG1QeqgHGBIaNUJMHCKXPqWY4Y+JVJU7FKVkExm1jOJGwskV
r5SF4j9uJbXYYs3ITf5dG/L1TVtrKuc0vayxQN+0zIcTQy9SY8rVA9PIHfxA2zvvbm3sT+gRQhmb
ZhEgU/rJ8bIb+aORDGI9RA0RPesRoCh+g0lAwDqXL8dxUFu9BJB/gEpT6FKAljvLiOpnC98NJ0iO
fqP1xZUS7CQBnDS4jYK2RBfScAwHphKxpj4YaxalSGWVW2/OZng5PGCDVyjIhgKw4axQMp5ZfZfh
a0aXA7vF40mO0gsK06PMvTe1kpECNBgcVejpIWRKrvFX8bSKuCLOTcSgAW4UGM/tdsINp9wD01P2
UMR2XdUKcNGWTA8cXpqdrjnbHx+T7rRfJ/oHTXGiQl1+MSAiVDTcs+Lb9O54n30v30jhGTzIHyBM
0df9Shp51hDcI23utRfWp36SJ14XylHbz8LgNNFghfvMv/8uMTA+PzWwkMjELgL3OEIxyafGteYK
em1TIGbFUlIVR9V2IwvpgPm6qZKvRrL3m60NY2uF5T+LR7aNqwssId3ZzlwHfk4HL6p9AvO5NNH5
rukwSw3H8qkWvfe/vdR1GiTXKF5jlbzXCviv85liMbHqBKBzeKZ2oD39oP/BLi0Doz6PPy24LKOY
x1fhGYX5xTI4F/+4wIhniswgJZlpSBTtemJfC7zi+UrxAtwkraQIHc6cufqSsyToMGf8tfUeE5Xb
hi6bVCmgRbQatG91NxpeG1glEend9zNyODNcy4ACfRws8ejaCfCdL9xioVqJjnAcEzBXVWsRCCwc
qoStw78PTD5BaM/Ypr3+iF68AVGatlyKmjfOGYbOm7tI2jLlylwIrZGNyGxHH2supzZSQzsF37Di
aYa7ED3lF0LPPlh/fWSgUbT6ChN86QeCxL67wASLG9yoZ8ne8Yo48oIpkiVMQXqZib7e281K7Qpo
lZQ4eB20hvq1lk7frBLV3A0hvHi1XWEVKPG4hKJ3Tp5JT/Wx35FxPL3Bv17QLv7NV+XOwMSU29hs
4M5LoAMyJmsDkhnx6gjD4p38hUdTEJAEuHDekLc8fTKEcYEssZQIl/Vw3cf+EwbGhEYujDK5XJiJ
IhxvGVXJ6XAQo6iKfiUqs6OhF8hfpAqgSJQLQChopj/1lKEMIatAWMljcRERgOenYZCjG3zjOgG3
71uC4CM/Y+JwlOKSYaHqV4Jr0hh+PmWF7sZuKBCLiO4wybrVEfmJogTNqu1NO3QnUXn8ZRI1cgqq
Lz8ahx23tNh+y3aTu7DD6dAUDaDIqWy9gzod4exA1Dmxd3X3MA4oeeqZ6Xs7fAefvqkiyUZQdBhT
3K2PQx27QcExU9bpVgieXVqmU+KlOHjYi2LgBlNl1JpbsPUamGyF6zL8XHbLmX5Jf7AA89R7cRWI
ROgS4lWIr2E53ZU16BeDsce1K0T6Fi4sYI0Gonl2Ek0wFjMQm52wInYNlnVIxSSb+7scVFHFairX
oLnTT7sgFJM0l8ggo+gEkjbRq99zn3rrM1nOv9z4g5YRifniFkUW+ObwrFg0zOjD+WBx+QLKwtbO
vvOHEnrvTW2ufMGPei3AIYfb0uQSp1TeMepp7YsHvyjquZNw3DGux6wrQKFSBZluol9NChijKHRW
Ie8Jk2fiT9ZmW+LalWKjJ+eQ+lbNtztswQN46n3KLPzDiVJ652ZJ+8AyAzhR4uxg+GFa3hWgj6ix
MmURDUT48GBzLMecV9pzo5/KvhrkUuV/y1byLVclajLaoGDaBsaw9TMKQ1hQrZF7DMicbL/t4Ygw
SCfMSsQv5IRe3p1eF01CS/vdVH/OJmH3Ud/KxljTi9n8UzJbqZmb/Airplp++NiIO6Dgpklk9cTo
E96/e1n88JtQn49654PWCp/WoV9Y/I6MdUe5a9L9agDf2NXn0D4JzV1uHq0ZdtvJBmtgOHHyw2p5
k6t7B5i1sSLYy0j0eMWAF82GRxdzLAY5wwnAd/DHhQgMqONmq8T0xQC8JDcUytedsDIsurzjeTCI
vnhqImLW9AkNiEIskV053XU/HP9X6GRaSOTDpnkm/qk+muHjAVWFHTFF2GgnPOp3BrXc+SQlCFBs
rOPhsE+0ZQtw57WuWbv92I1uYNK8nJBKHZqrb+4mi9FuboWMQ5kbSgG2nsLPEygxWen3LP9/RWu9
vRE/rO6Km9FmD/yWJZv1dkQLnkXibFMblVFRd185D/Jmv/8I9gQRj5GwliZcsDNMjeDVTxjPkyZB
M3d/310v3arZrVhi/7/Izao3k9mYEg9FQHyhLzKlCMSuAz/e6w0qlr3JBMvUUUt8iG5P5By31jtr
kbilgFF7GUPArCgu6bz3lzUulbXyl3FCY9Wx6zcbEMfS1f5Pm/SYrjHOtEQbvH1UvTKticl2koqa
i2nxKMqXWa0Xz1F3Gj9bWPSohTZS3yOhUbTQOz4pMN1xC84h13fmlJIXd0rRvIw1RnyEmakkxoJr
eus9OCPHRNzCdtjGDeFnS8pCuPFX/qj57c2w4lWOUqNOO4r0bWgydTEhA8ipeV0l67G+wSdAyq07
/ge/Z5e5m2Sg+qV5ON/3uebskdoJH8yiZneOIr826VwsrHQBVgk5e1XRlTWYEwmr8R7RMH+Ctu3a
zuV8/8n6H1CInWJLVRt5FAN9xYuss6Wy6plNH2uUWaROjir8V3Ez/ezyOGFqzAjs9DSFquHQSXXS
J7p1lMlxojMkRACI4ApX9DiH0iMcAtzgImfyw8021WC/Bd81caromgYaWgJqWWdQ7SPOELH+filH
ygP0aPf/ri8Pzn3jvKSzxPM/6VKLWD4rr/bznWlDCllWBfYKoHLxnKG19y6oxSEI0AuQb3FCvPJd
V9vzvS1uCpgt1CNuZ6qKdTs7n86fNrctvNmcW1ZIik/O5/thYzJlQ2HJSVTy63dR+40ZfTaFaEju
WjfvrNT4k7DA8ngO+BEsLKN3+DlCdNy3AEU6T15+DHwSMixeLfucz+ACwmOEuU7gL6ayFgxgTPYl
FHqIlM5Qd3LgYTHqNT6LnvP6vQirN8sEK6iOskWIiknKJXdes21szDQCw+GXX921lcPcNPrqnDO4
TB2pBFpDqO0uIfBbG2zNzSU48QZ6JLROzeX6jiwsXXJKAQleO6I6K+rvHsY1RRMoBc0M76d1q6we
oaCLWCQ4/2DaIWHIZomORbJeom/auVrx/6YQKrR82dCZ5cN+55EBfobgbg197tKmx11OSZ/immLr
BazQRB5OdUOyotqclaGmIGMnxrZUrxQ4iSUOhMCPrXTasfnLQm6+5MYHT3McqR68/O4Hj219ADss
zwNZ8N2/Y9qguxTxTM2fsDLIVJ/oIrxKRGbq16kQ0zCJEVWMpoWE7egelhnbN+f8LnWP6X2jvUze
5c6dukRLrivVSZ4/kHH4D61/mIpxDfOUSh76+GpiqapzJ9tRMe0It/dmEb0Q++ONWYnNZR1qyUFY
gRu0cMqCGSlZjIzO8vJZRH21zGmd2nqfRtbfpyn63lPRC4zIlYLf1zDw+YiMls153Gt7g4hHlObe
MrUeOSSjwt/AVKWWzfTNbfB8kDhqo4fRyb0D4UhQBxvljT4UVZ9W6xqG4oSDCNWGmh1ED+DqmXm2
35KmdiubZNtYF6cU0RtOwX5Dl/PksclQPPBSBC6uiAUTCYyvyplibNMfJGk/uPWimNlNNT2A4su5
Jyvlz/j8ywFBoHb8E1SGs/MY4LCaG8tvkC7+f+TPUbWZ+WoHkR3sRPO0t+/xGT3cfFFTwFvvdeza
Kppkzzpw2MWpoW1fhHCjbBOqZlr4zEv1g6HMY6JyuP+ab5Pkfl1DgUMwPzyN57MT2grsvdxe3SdT
rDOg87F639JqklppWw8BY6I/ITvIchNg015gWoGNRy6FxcAwD5Bmv0EM7HJKEORQ69Tgy8QEAG3g
K/EeLyWd6I+j0jP07i1bMargzm4BQC4V6m58/p2aX3B81za1ACXYWG08FgsQQN+HbGVZgkGhjPFR
03ssfgFgF08+gO+CWOYZuigKRiMPUuYQfHnh9kIydDlW8aIgW7E5qQuHUz4HUUIYq79xKuwXCyio
9QvkbKilhNMU8D0N5B5UKfmI5Jr05fLsdCdIw8ZJwjhLL4e6QqtTvgO+wc32mMBoch45e8WdG0GG
4u/C9J1c5p+9SVLIKSo2YBgTrQ0HA+L0pof9Z4Ju+tIp7Yankyfbh3Wz09DVaw19yy+5I99HocPA
y7awuKe4tocKIbl2OhqB/6+qC8us315nHBAIBvojNFU2VBgFF7xkvIExzJmJfgOSuSCuyLgeMsK4
N5Cv2ReLnlvXXVH1sI5z1SIGFjOBFAdQOYm7WDimtdP+UWVs61btubEX7nt0O+bqHTKfx59u4vd+
LEolIJT34Wi6k37CbO7my//NUJcQjLQixiUCVF5BYgaedI7ec5+PD9Mn0uGDPaZxr5qpLzhGVMe3
E1np+b8LVs/1trzbhxQs5lf7uXyDTCZlrq9AQXvMAOKqc9zSUCgLfhTUb/IAElYMZDk0F7/r+XmA
FIC3MXPyCMzDD+5qCMdE4U5jAe018fk8KxXB1a1e+/Q+j+A/p89VoA3HUcmLduDhD4Ckdk5BHUsj
pOpWzlcj7LyYcqAoD3pRluSID1SIP1KkcwnuugA9drK9Q2lLfsy8iVLI3ENuBYReTx6Ad3BsOTON
43yuKrWtO9wUy4FM8aXaEM36LQ7W4nd0N216OJfU7X9ULPUJchiFJ4nzpWhxqHhjoxQKlPQjd8Ax
M6vzrlR77bZYiwRR9XGDoSFOSKQzYznPNqsKph981bXzh1JE07jv3kv4SAyQzVJNVdVxIhv8VNZe
g021ZrTu3SNMcqLQA0/N/qSsJJ/GzriTX7uBVcnnDbIc/HZl9r5ufXJ87iYYLWAAtfqYcttZKE2d
6h4/jIH9eHf8HSxaHsENpMP9grCJ1+yNitQHCvhJA5fT9eayZo6iHSqnQN/D04Gxgdzx6vf7YdJ+
zZArcjhjur0K0YGgJRVz2q+GFKq9oNMjz2h12BnjTJSeIBHukGyut3kjL56husLI79Fue2ULFG3B
z+bVWXrsQyG73Rv2snMIHk22KFyht3hRJY4Bmi9G5PPDAU/7xm5zaLzpfZV6JF1AfaS8qAlGo6o4
MX4f9F4M3lxFCNgGTy8ZKDj2cLf6gvCvudWGT5nFmQBP9QlfyvCVhtVV6ID9PUOgIEovaAg3CsxX
Uoo9hmg4Ljpoplq2RaW+XmlABzWXCWwnIH8IPFXmkdr2gsJV8a89VpCkqPRexdL38zO+bOyf8QW3
bpMby/OlEZAiW16rrDAiBX4YrnIgUYWB3juXd8NSRyBkefGRyMBufLibz6uL+CMeZnjKF2j8r80e
snxbs5v4B+7kUNdSgqutj23MxRTcsb5r1nzpTcaus0PA6AnkRIjkP0ao0vq0WkejNpDNkwCXX26S
Mr4MpAJCbKqYu675+wRZmek2wLnXzrVudUZ0GeI9oeF0MfLo4DdjK/LbUfDJ0ARgn67cfec1VleI
X9qnCHbitaRMvkCd94o+rRgl188bu66Bj8q3OtgMB6e30SzJYBYneaP+eFad1VsAEX/Xqw0IZwjW
M8nK/+y6Jog+X1PuEuZYccxJElR+RgYztueHKTd/BLOqJr98jhKh7xGiPQQrhmQuxZktAjgwjX5t
WNIEUxCj/EzBUm35PRBuieH8OySHyTq4EuctvmgMgDZaT0oZz/2uTAA+EzCKhWdYaulFwuWRUADL
HcK0qU9UDOC/idhyEN1q5jJWymQs0PzgTc1JjfZnkDKLU8E5AW2XciJ+3E8mO+8XBbVH7UzfZ/iW
Uu0qryCDWgJQwgq3oHHXTL1JTVvrjVOBNu7nkeJZLqa6EYPyvRyYsCJdZKda7VqFfvmoEvGNaJ/y
LTvWn6Y5Nckoc7GL1M1LkQgxvMkHuRrXrqDMBPB5wWWb+y3u9Yw0/8MVwmSbGf5lE5NUcn6CZrXj
RCrLeGA3SJ0mKgqrFcvdf75quOWtb5pQg6+iiS6IzhzbLrGqmsijHtceum0kuTIzO7qKiFlLdnAG
8oOX/N+E+NRvatrZsUXhPSgp6eBSALi+CqklRKoQi9YDJB3hePkt9vAsow3I2ADX7Qhh/pkUyaxt
4orAxi7+qU98XTUFYlfm1GB/3GwTRZD20Hqj+l2ws6lBOHgbMpraPDnny6T4/QMgt51q3wi1bl5Y
0q/XZI25BWGUrQ68tN7LYrrhDnGk251qvMroBw5Ju0t26To51MftaX5q4MytYY1B1Vrxt45CfQT4
JoNP5G8IdhSgxc8H/MpuYf72tUOcgdUaJ8cos0jNjiHqVXnIFecq6gcASlqNLEucB6sP0petL/Ft
a4ovK2dR7ZIZXu/0rm5BXKj5dcGpVR323QO1fRt03JrneOMvs7Zth3Xw/RTwzWVhoegJcicJByW0
k0E+i+h4rXz8V6vSgP2OZ4Fi4XHIDyyBgVWqRqMNas85O4gqrgbp5C1noFGm43bHa3L1SMbeWBR2
5vAVl3H9S2PDnzgyQH9L+BiJIChBpUi9eKe76dxrMdxYUjDuDEC+pEf+NCHSH4f0xpN3QxZl9ZVJ
Vc4W7F/nUTaLU8Ajke16032zOnoChwWcNcDHkbsjCwTOkjoiez67WIx14xAGQvNscfQ4MRZIFfBH
UBG5hOdZpRrlfzNZtnnuJdmyExlNw4eWwk9D/AThSFQPgIvnIIuNngsvOJI2lR8MQfiulGJf1PRu
MugRpnWeCESJL5cqNHX4trnwnhkBdohQcXwiuJHQVTqPj54KR0jTevl5quNw8h689imAL9Xu7RtS
4MAuA05yuXfNfajvk53+yPSO+IrND/HQnjP5tBCmoRuNkwyy2iaSf9iQyZ9CUjfpMjR+cCi+WARY
qlxv5A2vtUmzvFhY38ZAMcXPJF4pPauJZ4xWzTU2W2iU9+szUo/2Z36fmaIOJR7YLeQpg4RtlAYq
y+4nJ/ZawMVvFK4igoH4SKQE2MMwwGVjP/8AusVhz7i6/BzcQQQrl9lnulpdiePtm2XvAPGz8c+8
UX6NG/9UzLls22fTj3mIth6LJCU6V/Obd1jjLo9gHzTAsqtMgeude/Pe4mPrCv/8MhreeO/4S8Wn
2xHDQAF1FmvYSRUW/Y6EXgQDHNb1mSkwZrs8CzCaaGAa15pTDAZ2ZbSe9VlQTE1X9geUqwqH45CG
+o0QETkvJNZ4HSxjYfl3jKvC83XhhB5qfRNddkoQ6JSEhssdFyxKZoTlQjuTXeFElcVUtaEyA94K
Mx3ACcRWcpNmVfCVkqppt0iaRayZU9q2bmNkd1L9Kgf6/WbaDmBkv8MOz1Y34x7qLbPbPuChOAe9
lVgnUPe8HbYGZc58QCgxx5lJBESl6YxN0BNxpDfNrpXsD8ST3Ya9PBoiXrgTiUo/zAuvgAmlqpx9
YrlX5wWyFmFFyYo2wSzK1LxSkcmCv5ivAxRTd+F7vTfjimPu8B2zWLXi17OHPPfZKNEgCamXUfN4
KACURgpmwVx8Pu+1qjYbY4I6GFAKeQluKRKX3MvLuXjcMeZKxgIPHY1VzbuLSacemz3GjULlv70C
hXVqdQV1VN/O2FVyaK560clUMdXladeZUEl1uDUN49FP+ao5qmEjkLB+sutgbEolvLpDp2+oLnbv
YzRgmWBW4yKaTqhZyDBX9BXozgW0BlQfdJc4uPGWUqB6gX07/BS+jZjSwSDrMwFfEkwKkc4+cet1
xNmDkP+2lyVcoi8YHVwag/ssGR5ULIFbwticVunNAYSm8Lic3CF3RVe4ji2kRARmhPBLNrnbT8yz
pzCrL1ozDH8Ggnao+s6TsvesD9rNYoFVRsU6rtKXQpJDqBh+Fst4Gx59zWg6vKu2IJE9xu6hpV/3
5M6QjhNHtRhqefTlMZgp+bmUXE1+ImvpjMkgQinPO24fcThTHfLbN2EsXKUASssJ6UE64SiY8tF7
O/GIO8J4pTyG4PVLJ9+4d7KvGclyS3y31SwCDqnE9nK3B9Vza1ejsNNHCoQ9lljT6FNLKkz17Kvi
PxfJMfgkgupW74gRQHgkx0sWZ1A+Q0I9XR7C+H7fRdbvwP63VktThsg/39tjAkSZOhINZ6ZVcFW+
T2eJ/O72Y4J84Ac9spqSE+wX4sV7omEQbHP5mC7UkjEgagKNJGOK6pfO9fHh3qQB6xh3YalNEt56
9ARbquZEC7AyK3oE1SG+PELMA6es6DGl42t9JXWHygpPyuJ2v7tPox9cvSg44I8MW/X7xqTD5WbR
7a30wUsgHNY1abw0V2JRtneDtQLs6ZxJuXyA/3HE6LCuAx4DOoZw1oU40Cv2uw3TIzYzHTJqC3VU
2b2Ox31vV0/0YCD7eYFS8kNfXLq+t+F+dEQp9c80iIWJzTjQYXPXexsSPr81H+tguudVqZWIfdJf
khMZ+Svn+zJe/vkmeVxYoLlGOxiyJYqezkL7rgtcgvmjysgXe5T+N1vLxuFg6yRo2J91VLTSCArx
33um0b2hD5kXfM9/xrEC1H82yDrTiuAvPIzXqmzhhCwU5kUiNaMa6RtK1YRfbLUfyATEvPvElKW5
G1rN1F9Ff6uWS6zlLwLbgWfdmDkH090A3r1DN3hNh221BiEE+AYpQkZ153oZIaeSJx3i6MKuZOTS
I6zQa2XyT1IqjpJaRlspSlvERigt6utieCuPnvQGz7JivQnAd4UEpwjoF4m5ixXD8Of1PhRy6CnE
v2fj+JBNEJaiJ25f0oPjc4T7ojk0lIEF/8Ac5ru+KfFDEhWUSzPh1T8GeXFhX4s3ZLIeQSmtw7Lk
JCj/AGPrQFHXhVXTVjcIiVaKRV+pVufkNQmPff5pY/rgW4XHumD/cU2ZMGDxrm5PfWulMiNqZt6A
a4e6eHYGCUAxg1xl0RMK20HrgZuwCeJolF2ff4+IqCnISQbAE064KbHY8shmRY3LEe52gCWQPp9I
f41ENnoU039MN7BJlMqtIYt4q3lhPMt/3xbAakm3ONy5i3NNbR/8whudJvv7TwETQ4WaAXkm1+pJ
Bk/2H6Lzkoaf6YL2iI0sfrtEgGc9qQv5tGgzSbe2xSQo1qEBzfUFhSLtBf/hLL9kxrqklaVHGJLK
8JtzfXuw6nFCVSzgudC5BVhra8k+EpE6mkQUvicPD2UIjcVZ08rtA4U2juSvdkd23iVnBy/svoIg
zmBeW37WcPx481LQ1cFrfvc2aY3AmFuT+Fqm1c4gTcQYdx1fZKZKAKqlHWjs5/FT9MaF373n/Wsi
iuJxCtK4BcTeEyzdBshDEKPRcT7NArO1HTLD9IMK3lNZMSQAjOTkvkPaN5mvW92muu0YflATCiq1
Ivio7OndmOsgD4T8zEOiiiBejv0BS+XS/F+FiTZKJkwnLuN6UDSMO0D84J6YRilqtX+PwaByBTGC
8lyHwV2mMOJrTFeqU43tY3ujz2B/hFf/G/LG3GkEvKwfPYFm2QEumu0wUExG+cJiXakaVgZb+5q+
5AGfMKguWlG//tW5bviEcKTRnZJOZNxPvSMXZvpEt4oPN16BldOL5XmnJfTiBlomkWape68FtkLn
dH5cYKgVEhqjx4J6x+/NFtbUiPK9+kU+Pf1SKIrqUfiH5K7jrYb0YEROZSKBLRfUj6PxJ0l4OMKD
NQfhrUjDvO02yWRa+hPmjdy/i9mwlNiJXJ2AoqCEuqsPDAGIcVBGQXZc6vYzU4qYFLIRQb4QKj8+
lj5kTQzTFImjvc82W8qaiPpW6FLg0P+v4vAWNRKJKVv4jWlKNpckqkYbOxeM/2RfWqJxhcsq1q+n
iq6nkBSZ9G5pFKZDBrW4Jx9R7bpaccfnbgzFg8JT3EjLuGprABv8qzuB+A6e+i4h25P2ywv8jnbu
ThXMXAZmJ+sZXf78lUx5XD0xjs8Zt63sLzUgeDAFpEpQlfhMlN4M3LVW/XmjfikZS1PISRRaI3M2
y7Q64OCOBaWpKpiWLwVyuqvF5KqnnfgI7uUdxIQ3qds7C8PaQnkUdiUaRSpV3WUTMjze1Ta4Er98
ZumWN13n4qjwIr5vBQGWgPO0j1yyGwTehfzEomnDrUvVEhgLx2Ug3giT8YCSIT8pWNOWgoj9Gl4u
uUBV9UGwHYnSn91ODQseriHgyWpoj09HMncjUAQ6PdO3jNsK1+f6zsgAuQViTsUqLRbatO6/ZPNv
vAVZQ+ZiVbQ41NAN4yzrVGOM5K3FC5xnN1DVwJgapSxR9tL64ImcC0Unkrme/qYZvGszSa/f0DE5
niAaTFLdAspZ8NOFWj13Ri8sJBPmKDu4ciXwvkllSaRZU+c65Piw98EGSSloY6JvOd+AOq3Jetxq
4e4EjqlGE/dT2P0QYotTuF0PAVY0uxuvLFEG3VTea6g+SJB6+H2+DAnxttLsdz8BtbyN25dZ2Tvs
Bc1/IvD3QNjAg0KeA4DT2xfo4pWcg+SPNxm3dveNEx2TA3nkzfuGEv3KH7NTZA0luxmDevZHYMMZ
IiH+gKUg5/z26RzofibdC89d0SLFkDMyZ6aeAjo/8j8ESiLy5Z/LosEfvpcmBpA8eANWBakUwNvr
p9pbw65/69IZUBXO9xevbkzruru/5XsD1s3e4CjktW1dmbOd2QuvKCDEjJIH2ICCYgAy0QTYRXOt
nIPtIS7ULwHIxzZNp104SpB9lqLsBg/5zvWaFUf9/bMFOGwmjbm10fs3bJwlYjay6L/3H8EV+xV3
izVMjxhOVY5ZkfHZYux6jkWDifPjpIkv7hoRUyL64pRfvaH3sSUNeXQF/G7FpSUxOBg6zPPuX1ze
O0RN3tBB49BPk48lfwIswhed0r7w+9uTbOiYMX+Xewp73h6ho/lnuGmBi+4tV8ANNi4vI9c0VTx5
q93Vve+OhdJfHRCLSkJt5Xx4lNboOoYR3VML2rBhyCug6ha23MZT6+Hw1mKtMOVmdPj0ey5LhxZn
E1AQ6d+88EcnxbusOoSuUGTV0PTJ3vrZeVBEmb4eMzSynN+CH802YsO1YrLqYVvb3FC6+HEUGiOe
qweApzxZk6/HUM9vloMh99Zrt7+sChwQ1Hu2uh8YYYz1Gg8ywTatzaCvC/8uHZ59XacGrjpW+5uz
Sch0UBJtLtiE73XImQC0Iq0Ie+VZs/t5zSRJ3urWXDnpv14Lew8zubS1/zhRWGdLz9Q5pZHO4Gku
e4PbgUiSrx40SnQI/AlC2ZOzwic5K0k8Qcwpiog62vTRjByAozOsV3ND3CBFmy39B9wA0UyMvafQ
1pFqoPG4My+mjrHExYCOKKIDDXdN/9+2YzcJ29Pni1sK2zjNrxQ8CKjBkFcQBUJn2O1vNlzrP0tB
TW2AAI+LVkVIlO8/TcAUc96rkjHicGo3KOqQcEcTD1Zg/SqnSgngdUnjrCaL5qGLfHdDHCp+4jDZ
zWiuW5OK7ahUrUPSEJMIefJfXEHB1IUOSh//ASVt5Ny1FJRuGM6MU9DMXXjqYAvow82uOenld4e5
CfxP/Wt51yu4cmr2UWw41pt5/W03fBZ5u4zC2PBjgeOlzocSXdA+QFFK4vmviMHDzYlUh8t3/l/D
P0kuTm0NhP8L/yoOegXQFLSb3rl7lMZFxrbHBmsRjFUx2djR1tZsT2PpuzVfll+Ey0+AP/lmgBZE
Hbv3LJBuha+J4qhKhAcYNBoC7lgeGMzrhPzoRHkL7B2XwxNgL6hZq5oivSjgrr6LFBh9NAJRJ0AI
njbb7qhOlz+6Vn8ZG1iRN8ATV4ctHF4zXOcO1N47OagS+XyrKXMvpxn8dUBBqaP/Zs8FuaWS77gf
Yrdd3wycJC4gMS00giaeYDsuGSV9cqvhy8VPk2y9hnC5jFSSzdZAEgvKYRtJtUiGNaFzMcqecgR7
qxEIQ8pX/q1lDRRd8XMyR4LdZJ7EoXb6BCGsle9tXpXA+VL6OJerbR9MATqzr7PeiHEvrJXoLAF1
XeiNay/rZ5/boZf1jvy/JQ8oIktbhJ8Vme4t4DsAy6dLiokG9A6+jMR8AvZem2XOiLpQLYITnR+s
Gc3BvTMGjOE5t4RcIXH1Q2vP37/9PZpylXdaAaVLCi2WaDflP3kyv+kEjDyaxA3RUkCfV37Pc5XY
l+ENLiheUC2hQFFKgUqnpoU85Hdk6ppHbF9Kpsqc3veeAz+K6V9WqnSQBiaCCon34UVsTLvn+L/N
jwrU85E1459kAh21hmU2vzLWCWoHm4WvOAmDmfdPoIcxmjKgXC7Dph3RGEzZ9+HxeuHqxGLKIxXA
c3uD3tWWUkvD7CHI5aSEIa93V5NQRJ/XOKe3juUCZU4AAiFyCfOqVZwubYI3XlCRLP7AeJtDhfki
FQyIDbJpHHN24G5jJXvV0aAFl7ElpAD+WNFEaCChxj4zeY+1OyHqYSCHmycCFSoqrSk6QDLxkjoY
xRO+potnUIGVnFuytbF84N7Bz1UP1Oyx6Xyf8Te0iPRULN4VhdQBuJ5wMvv6DmVoM6sLMXXlGXJc
LINCl6EKLQOsYf0oeXPU7lg6qECCOWfS4Z1Gx0YHSn1vmhIAFpzybOGIOnN8XXQEVA9p2gxEXwGd
iBR+ws/vFC8jlaXBdNOcj77cgZtE8TnEWP+yK9R53XMh6UjY8gi7kCWcJilUV11l5RTBYO8LkbIw
hBDa/0fpSJyFM3LLovtFn6wKLEtVzmmPgap6RIKzWSodXH/J7Dq3BN9J4TUyusZO6WWY4fPKO/Yn
u+6T699wiZ2JcX5MEMZQwBChuqxgf7yUbN7TsIzlGSFtnqA448vdbDA6xRpcCCarl6JxZgxoad3/
7IZRo2ruU8laJo/s1lzHI/EPe4fi/UCSfATVCcHvyUEw1Ri1B7EIJjLUWtlPWZhMlVWNp9h47Wat
s8Iw7NVo2r6Funf12+w2dAkegpXpfrdDep4I6NaxgxHEIhfNYDhbw+9MY5wr8wfNMR9BbtIu8qps
4HaG5kX93rteMFJgRmkb/bLSmftOI4rV2+hSEYhUaOrQ8rmD2VNLWWUXflanA4E0dK8y2Sob1vIV
/XPIS4y2bKbBPjqcQwe/A0Ke9Kh+qEckeyoyQza/EdWATbJTdbmQ9R/6hD8fH1Q+fFSyCkSrHXQ6
WySsJZerTVkDtneDJnHSek7OzWDThjtO1zuMzM4sFOwvmbhgODwbC8DcxoAYBi/FVje6dtpghX2k
0rL+15HOcEVHbKv/cCbhjn6552fjew9KGMh2OX/ibzvT4ZAmp9ksVhiQI8SN0wnnUXJNcN+WTWlM
X3Wu2zfbkakMp0irtSVvTt8ZHn0h8bYQ6fVfGS4MsZgZLUrQ8/vEGq/xoFVcnE2kGPmXty0z+gYS
pkVLPjrVvvwwZTd/CO0NeaWZps8+rvQ7b984GLGR7RkDPkc2GJRk6Bj6V3MvwY+EemxQ8chnRo+j
TmPgVj/Y2+4NHBq79R6xrTX+O3xy8SmodZ3P+KcFq2KKSYBrWfv2BiFHBum1q9ZF8dZaG8bJRqKo
cI2dNZ4B8C6wHhe9aF/zeQg5N4DSilXqfhxXIdj2sCLApX7bkMtTPBa7c4QsqXBg1OW9BtWnOl+I
MK4Ue78Utmy+fZp6vzhIvgyF0L9eTu1rT4ENS4FgCIfI/C0uQW3UC7TmIptQiva7ZcZoxwfaxm+u
9Yc6Xgjz9VgBuAvWO20PM4uXUrU8P0xvUIdcEYIjHM+WBvkHRs3XDtkbLaj4DtDnQ3GhXgIUx2oG
Qk1BtIo2uHhB96+e4FRMyzHfiFz7QwQEw8Q9gDd6zSbRoKTAvrqKOf+kipbYORn3caN+WaiWPSB0
hIMRCyg5waSEckGVO5D/krTBVe603/gq9Gn4z452GheM6EYX5DXMMkHJ8qQtdbd+GTtVRmagIMfU
RHi/MCjGFJlPyVqgMAPoeTiHa9RUzAdPgULiVQ3UF/DQttQ/xsEIa8q7xLnarnjTf5tZwYmHCIfv
E9FgNSkLiirY4NSr3XwMe3foJtSO6ueIkH8/tlCnHR6z+UBNyY1w9wgLTZlToKvtJufP4QkAYu9n
cLEZBo412duF4wxWApO2KLvqhFWemeCCIYqrYLc3yEtggJeOySM4EdyxQB689NSQ/cNfHZ52GIYD
6vAQUqhU+kzw4WXbtP+9hJJ8tUtHH3d+xTgh8BegLAvpLfJWLm1X7YaEDbsbeXo/p77vbCLUF2bG
YaxSUxMmKqJrRTpWk3tj4NV//k41CVk02CZ/onfzrFBJ2cL+boDAHFjjnuqCQSZDvzHAvLmGPtLy
e/6WxiDJuwKl9B1WorkZ+ebXZoLpuWtz9qsAETiTvupA75Ea2hvg5x08r0WNQI5c4r6odc5QGyY7
UFXQyTxLBECqoQqDkKLQjStwbioC4/AzkCBv2reqD1CjtPlr9/Pe4nBgIxXTb5r+/gWv2SITxs2R
eOUopNfAlXqxYkzVS4yMMIG8K4feiXm9zcSgZBhIBBrqYSBs6ldRWQbQ4g926ygFpmzqg0/L5cTj
AsUHmZUbhBxIFKHxVkMYQYL+Mad7HtdBYLoJSKBGbF7XV/vWM0b8lsr76Rg7gdyVlx9sAqribiq7
Mu+3dRaGNYLrIHG4miXd4yIEy1VqG4VLKpyJmf8mF7OGl7fwjxXfkShIIQciSU7Y/oy7zL7gunmy
wCjmYKFj6UNxe24dU8nmEfKZEtqgYDJMHKzQbOmwypwjqHhxIWgbCa/59/6Om0DX5tWlWD6MoY54
NCj2P8kHJq1sbZ2lp+kf/VoWiAhM5nOn+7CZmIPT631RtrV+syaKcDIMbXQRDrAm4UzunIsyz402
pu3H1bM6icG0ss87uLYaxAQ15k0HSjamn49sxP5p5N4brm71wGFDsxhE92S82/dfKB6nOj2wy4o/
7NbRcVUPT8Q10TXSuToqSqtrW7IqzTGvmy8h7+tU6fh0rVGeUCPKOimSi97koQJ0om0oQsss8TI2
9INDgBhAPYlK0MbqVMECIPoRT9rmed+cnz23O+S/GJP+osEcgFpdRwNrmLPHiK+qwzOL+Lbc3q2E
w55dFIwBFU8opHkqwTiho6oI162X+TLseAsZzEUm1nBC4CvRO5mQlx9g9ifuvVkrH43Kd7MJ3hUI
uzDQuNi//o+k7ljWVFikQHWGPYIlg5qVrSEQz0NO7TT7loiG6lcxPCX5YXo+REEmGuhzlVtmuFVY
O3bxiU304OC/hBJUC+y/y1xXsTKjiLSVFuGPdIXuAwIsAwUT5UwAQ+nAuSQh7QSPtn+WrDpz803+
BXBz+iC9ZThb57bokUniPKpRgWPttObbqKnCk9WrLeDdJXOFDetBB7nV/uFzkkWt+b2QHzY1QF9Y
CBrh/8i9DVn6feCc2piRrGBCGIcyzGrD4jF2oEfwCgwDoT0jcTAYSTNBqGCgUzRfWB1lQjPjicsR
leGgnIblyL1kimgeJrdrz15h5fiS0zA8aSW5KzhuPa0mxjyW7am+woRNWTm5J2JlS+c1vk8co1j0
UVA10QKxwVAVKKxkdbYnh7KFs4J9jfnZwL64qUpSyVaSLBfVxjL8MeE8SZ5gkHkoPVlqydaWiEwI
CMRfXYfNf6EPVkOVLD+8M/eFX977l4kW5uDGQhupmpE9Z+KqsCQf/q1SWLR2VEP2B12T/9OFdg11
uuA/R1mDCwB9OGp4xayTpUUalr8/SZ3wMDNgyZuZz8Tke7xewi2Kl8uN2uo5mgHTEDzUZB3o1VKk
1pmC7YCFegmZiXdT1zX9XsgeIgnvlKflKj7AYqAw0rLDF+D1E7H2ZZ2G2+SwVX03Ef55eS2/vOgh
beSaF+FO8NSkCgc92EliG8Y/JzwyRkAkyy8VagC2lPpMw6dPnN2eePtvBlG8pwKScDHYg5quy2yK
rNx3E2lrG43zOj4azOMPQPrXtJxGQeU/v2H3qX5OSxGFIJ/ltE00KzvIqRzrbNkMSuuZcDmQzJ8L
zR+P9Y6X0V7HlvSaifIlgFfukooJAMpTnpWRaXdZzHuaLOOdH8guMUM4bxHFL64TWgxKf3bw0fF+
t7IPMns7U0uy6NkiFFx9IjwKR8OP3HWk804/e3Vde2rPxotIF8mqKVhM59X/3jy2Ts6CeYvOCYlh
3b8n4YQNAhFAIXQzaQLEMYIaXNJW0Lqufi+OiDaqncPtDnnGqmdGIXTyin79sQJYvv0pJ/xmd/x0
XhxP+2HfjXzNDyxNWkz7T70p6Ml1NUf25GbMu41dZeM47I8GMUHsXER6TrWTszf2NsGC1im/k0by
6LVbCO5udifEiO8yW4+wRTEeemExegWJ4CGiuhPZ52xf0JmDyNKuMhi8fLozRS+DPZXpFepCibj0
YoMPMNyQdB5cnNse04Ra+3elUf+KaYNqHzR/TdTR82JZYUd7LpMK3nXopXRnXF1z8te/j4WSrTxd
L6ap7qQboiecErTP4jmZumyO3B8ETZU0WPCTYULSkIgVpK7natM2sq1LSyKM8wdMxzDGGN5VNvC+
gxWVGPc+NRdj0T87fpCU9G4qHZfTA2IsMJRRziOYq9jDZ/+AFN90eOuSgKv/mVlETbKhIV9UW2b1
jow83SXc4lCu0PglMNoz4ungJJrAQxabfyIi3OAGOAnZkqYKnX9oDKO9CYBsZP8PqyAsIxqXYON6
EeCEB7fv9m+jCp1qX06VPy+EQnugnORAPfccLH1LjVOLCKeW6A/aqdF/Beb1e3hrpj4PA5vB+6Px
Btak/Nwf7UYqOkxkJ/2BB6cEzJXStjzC5FIfYh09EqjT3hcLZevhhSQsfpmPnt7AVZ+odXA7oKGN
W6KpJvWCK3KTi6I5qS/oI0U42JLOYuRPCimk2/t8DS1Pcq5av+rBreYu8igj5GNcD+jWKAaKqVG1
LfVgMUssddayl9HNMJIlyEpbPYxYKFkAuODzYDBDHBw+sdXwyqiUY8AOyQXvOHlcVoCSs8K2gLuD
2nyZ0/NdJl4ar92bme3JLTo4rY70yRMgymyROHH9W0L/q2x8ITrs76v0iZKAG/XbuwTofOCmdFY0
rb9YncqyDYo1M9rDup47Lknsbv0wI777m+BCil961AyqCFdeyWoCjgIlKu3h1bLyXFZ9FQPy2OHl
3RzqK4d92PnEPNYywb8EPL49ah828sYPKx5xwBG89aT7VnArAipfk8zqPtpv+dIdVka9zlg7eQ64
C/EeWO7nE/zpbwjD0dN95el3CaPxLW+MkrAcJL5ZJr0Qm5kZUNptd0xhfUM2eel6oSlCl1KimBbm
VlUUbPF9BDOGX8dkblOOfRtcubKAPTBQOMElyXkSJKibLI6UCQpAkt+aGf/3Ni1b9ISPVMCl/pIR
Ark2JcWGspUIg05YqWRAp91n1KrVHOqxHhfwiLQxXfFJ7uSvpOG4tGjiVw9SnEUj0AoHQ/1+OF5I
WLPGeCGgY+0AbolftZuf8lxvipnlnzLGVEokEF0dEUjwDTfzi0uquDJJxQNZQ6LhUK/b9F1kZYdc
/vNWr+bFGUgkkBdKWMgFYzHxut2h/IHFKSZLFDboMmtogoVegMf4sVr6eZDOGaHfMLM746xTgDow
g6CCpo91eNAO6aocs1zzPGOHDu6p6j9lifgP/xnfvG97xm38a2cdeu2wiYQoFFG0NWfRAP8ITTo0
O+/Do2yV7YKckpRF7sZZwDpJuLcvJmea4Il8CeiMvn9iAPedWf8dpEtkRAfDsj4/vgNa7hWP3sPa
8IbyP9lG2FTzZGY1bxguwvtTdey5Gwf9F2IdxBtwVx1tI3eZUZOSui/QvdK26gH8jv3jvPg3gKny
NqNbGJaax3HmU65uUjGibzBe93Lli5sTzkjPrBPZJ3iRL1swhmAgxPqtQDcs4ahsp3ZhHHt0Hsqh
GEta63aEcTqq75DuCw540q0J2IrW02QhxCDWVLypfczHg6WnQBJBO/ef5D4J4R/6p8X+JeXDAhUa
IVjshWvo4sj7RuhOjacW0SNkJ1vgIkMOyuiYNXuORMCwsJ2jWlGQzn9f30ZFeeDWUnMNikdXjMrC
oQJGxgDpkIqpI/wnmZH/STJbsA0F69URp6nF/gt4t1ldreQl/VI9rzFK9mHowXoA0LI9gMB97iOA
eP0oAmh7p+9oM757vItCkN8bJUK0WcFD+Yf5Q8/3ZrEru2sP8IxX5pvMedHPgcfVB7+d+uC2LyIi
woLoSSo8+jIyWKvnO/ztmS+Q27xOrmn9YjybGQy56MY04J7oMNZmRrtj0bjoYU8J4uzA79Ke57Yb
SOtT3SRNEXBHRpyvbCkdBu4UXdyjEX+PcTP1WxHR9J4SvxEm5WAcyPolhOk3BSrTJMkhRxHwG0FT
uHBJsjGAbvdJ/TKgUfLM4PS/eacYOgm8ZihYt3t3X0DwnnogNYecxV8boBPRT7J49unGzRnaE+of
OIwVx4kRpdC68tTjz6VpmkXP6y3sh12xoDWUnVX2AuXMw3VBkdodnuyg9nvRj9XPMGq7wdubaN48
pD8+rGXwOoENRIMHTeWQP3ejWP6bXdICuZni/29TNg7CUQZTvuq+ObCXsffpwxuCNaojSuBJTPUb
46LwK/CXJiHXL8yGLSo92Jh1CRVDGOPgTZBvBbFEXXNDGnUFGyTv17ND815AtdGB7IOiaJFhyhjm
lJTOUaH9CtihkCe7zWuHAtnl2gsv3Uy7p5eXHuO4QCrr82ehB+KoBwmtfz8B/povQijJ9Thx1H1F
WARlZPjXJ2lDJWnp7lV9X086TtlsBPTFpl5WXPknNBdeohfbzu2z+JJCocZ0aqcUP98jbnzLTCh2
q7XIs7A+hwuqrhwvYyl4wS5ncp9bwbMIK305em8n8V5S/u6lARnMCoBpPld5DbSYCG2EFac9V2JJ
qs5yB4k3bJD6OBvYtLFR1HlQDdxEMM9+FPczlEWtFnfkssxADf7BXxSvKKvABUHPt6g9BBVZU4ao
IFShXc4g/hzo/d5E79gMIGWg1DPxq0B0NESAJGEw9ELk2NNJfeAaAhuiiMS9rDSEqg2x+mtshqnA
HbrL95IYhMKeSAjMNXbmPr4G/c89/v6JNjAoo0Il2NPdFJrBRFb76s3s372OtIlVkXvcpRpVxL0d
dfEuwNR+15LTFuPXPB9AUwV/nIsXJSaKLBwzv23QU3J1rnC37fEOAJ6TV/FMb94e/tIFlhG11J5l
1WXdftbIBIKOTKoLQRarfstEcBOz5ONKsacK9FKfWq7u44qvR6ipHSiRgji6SUGfr+izvSICJNf8
0oPITzecZpmWEubgWNpSXxPvrBxu+h5Ev8OZwX018PT65CmpL/L7mF5xQrpUdk6O9ZlZbZCDvagD
5KW5T5nVoPCJ6bUieFdVYPBaiD9P6QeaRLsvfHJdh54C4nI8xoGsVPXHe9ES14sQM8Swz0Y6f8FR
wm5Nftdsw3OhtklPQG3awaR5qFWDCN7DCRCwn83FWkP/uXh6UVRm3WVZRY49Mkr3sJ9qSTjOqcH/
cXnKGR9DJsg/NZtLqw1vpPYL/L9MQ+i7m8yEcVuXpQ0YJAGSJ+cfyGhmBeCIoDEZOzM0ZwFdxKoe
/hwhBDiqFYwXH/u5OItiOKEqQm8PDKfB+K7mwPubJ552pwes7/xxK8OB8jx7hbUHmb3cV3Xl200u
2YWWhXna8KADo5RR++jf0X3yGhfXsbu7nZiWOa+aZe2dBRAAW2nBh5fjpuBRbZ6Vm8Qk3dwBPC4r
x5mzLsx6PypTZlGEyCcrnd5MW+xG+baUpiq/m++2EoDRf+hVSL2ZhGyRNRqKls3Aw6Z9mdizbv92
VeNGRxqjWhlUwWMFfCMfIZMPUoy9FmNdhWmbzifmRP/NYNEtjEx2rC6VsY0UlpWTYzc6YzRD7Sco
ke4JCcybxQI9XhuNnFvMjw4t/7Mv71SIBoMz6gD94Fg2OovFpFJvHe0Fs3rEtjvgL3LlfsRDaqpn
iLY1AlecOt8wE/oMT4dHCVjQEI/APGFEe3oUy1jb+P92V7ONToHdPqeeuchxVyCBu7pphotIJVsz
PAyuZcUMdLvfJruf33psLuuVekKnN+555zWCQL4qXTMH8Zvz750Er5aRNtWSVaVdtObuOqyJffHo
fdD6xfQOm6BkgG3A6yXk6lFWdwPhTc2o6Gp+ZspU8KsXOl247SRxWe3Qzy1d/5tGwhxu+dn9JoPA
oFmZ/M9OZt9TXkQrWL51sAeSiQWC4Ntspmu3lkgEdcAvmQVJ9IevbMAOf1oJ/pZaSE6HxzOJ0kiz
e3JQCDUnKYUyww2jGRSLmft6L2i1cUk3K/mDB3kY3BcNQB+fVducxeFvBQ9nOUhtXWltR1OBrAA9
3lua8P2VzfTjkAUE1bhxKnK8UZ9W+ugBOgazW83XjapDU/nBan7iDcaLc/wOb5s+1vgF6CgA+M/3
JR4Qfqij0xhAbqTo12XsnQFJ+WV/rDcYfWTm1PBI7wToFANBsf2YjntQxsI9RHf1zs+rGGATDqTD
OquK/RNLQ6KfII8uVVg/Er1fgY8jP7bvH9P95NGg3UIGohn/He+y/1PDnJaeKhnCzyy+itxE63bT
L4oKMvAKyk3l32uxFTTWYnNumSIhEeNX833+y08MKMkCzogFIZ6msMxFBtSi+lyJ522xX4lDUVQA
u4fZyhy/wcL9wZ1wESsIpU5LooVKMF73lTVa7iZW3by3LhU5RSkFGWAeUNBuIpLSOChO0s7L3RNv
ymnAUIGdl/zcyl7J3W9RIA9ZnlDHu5HcmQ4nnLHKUqqColSk4l6oBNPMtR1h1O8OQfbw0RAXKQ7m
BqAzpuDlxLkn9+hK4wBM7FmiecPr1f3ZEleEfneElH/9Ymj2eVbJQAjaRAAowgKaVQ9IMyFOD5B6
Rd3dxrwqUa1dfm/E7UEwCBtK02z4VQgtmC6d+XpcKP/6blKX+7OkS9x0N2vEn8Z/oyiYmNQidP8h
R6OQiAhPAOS+chfejks7xFXqC6OF4IxSK81wtxHGFNfbgh4MUBrUsiW8gmIfM4RCu91NgDyKjIDU
X0T6f3xEYRVCpkZfTSvO+O0Z0mvK4Eh6Lh0n/fwCG49ppeLKKT14v+aSapaaHL3zsLJmOZR55aDk
ThQdCzVKXnFbRV34pa/atP6ZQvixO6VIoZbGpc+f99EYBQV1zjePMLOx37dZSjETd/8X9DlznBpL
Vk0CJKKpwJ76OljlAFx7D1M/xUnPuoAfL2Row9gMW7SU01rv0N0ii4At35GsA95CbzpivyiaXoLW
YSfWlpMSW6s4AaQtxO05HIdRHPw1dT/3wYjBj7Wu5Mr3wHkQ4IqYyAw+fnw11Bg5JiTuESND1D9U
HpeHihE2WeyUp69o9jGOwHauKJrko6GVDxJG/8pYaT+Y1ISVG8H4H2jadYVwJfHCKGTSwuXSR9RZ
8D72eYZ8mEmPoJ5s6Hh1qi6WBMEvvE603LpW3zeYcJOc8uSOMpxrtaNNRfoBHy+k1DIr+10TtfYT
hq1+yfMQFhFdgQ+YRhi/zm+9duIg00ryYjmt6/VyJO7emDjzinxSJpH+Bv5h8C5m1RBbWZxg8+8Z
XnmqNhNOtWhRImDkquiu647QWRwgWKMQvaYinT4jevM9QbWpjI4XjmcgztwwLpxIYOmWinWknIPn
z5PGG3FYBfD4qxAyHG/Q7j8Lyb4NCsp+aWzu2xNclqQ4dI2Rkue+IHkNrH0o02uJudDKWaMQSXOU
2tYrGZdyIXfBFV7NsPofinab2MhD3Zli5WzARe7YAOSusrB0hcberVx51zQgCEj+GxB0rO6tot+U
1zK/M5TjtWydO9jH+GQbMKeZ7dH9EDXI/GwmedUSDVWf0y8OhiSA61keedp1+Z4cUttExokkjaJu
SXtKeD1A55H2WURwqLsWvpIQJPeB2gkuHPZychlHMWcp9aIP6tXtjCE7p88g4pfeuXQ2t2MhedGu
nNyRbyIYhwZ3MCdnGZvQYpDS9KcFIQHvQEkCTJPev9ksq0JA5PnMhHxhEC06fDUCWLeMhfUqchUJ
x+QNONxcHoT5SIZopi+VvG++/glzzYY7ilu0JBPpWDZJOmP+aZzz6QZOQeq9AiupAFJpb+Mqp6Ib
yngJg5k/+Ds6ytggTEPmQ5ffXlx8dUcrJyIy/nlTzX0Xv2oPx2SWcEzLcKYfzLxXwWaqagHXiPZA
L1LneYrDcKMJuVDP0kW2eykKT/8e9i1envCsx7h9p46zp5CI4tf0fihfHe0b0dbPrUyDgdRHMEox
leTll3gQPpX7AGto5O+Fa4W7HWQ3oFYJQ/6PiasfiOsHqT6xKZdi/jYkukblbo1Vckv0lNXU2E2T
JviWt1jJ/MkaagfGCjGL7mJUnd2q9V/yslKCVl1E03iCsIyPJDQJz8bh6tLDxz0NrghMftYPIaok
pkzFw2xXv2HDca4YpYiMmaix2HtCAPwNzcvIStWXCicdGg6S/J/IuVsmUFcWRQYWuMwvma3ps90V
8JxXfthz1dzssu+j060bvsRH9yuiEQK+uQSghEsurR0zkC/ACF50gHKunULNWjAt8j5530b4o1SW
Nt7vIYB6kXKpAi1veeq+XgMbVDUm0raiT4VoTg5YE8I4mCtjaa0o9whOW/XXi43l2v2Yp8kQbvYz
UpbnRxM8Qiz3fzDKtHj3EH5Sg71EPXxkBjRQM0ShlxuUifSqYxanmwMNsoIrxaQybc8j8kBt3bDA
bgUclvXldBJ0BkUu193QtDz78i2GOvK83AWTGxTKLxHmMnGsNBuRyb+eUcTuyvd/ZD+AHDyio/9c
JXQE5tFZdShdKXMe93UjxaSBc7A0d8S5QNmLz2rzzu0fRXMjNmR1sBmqIUfRNeTHy7yg7h+V9Sl9
SJj0sIMDSTNNNmvzLWLfZxlMk0Tze1GTTi63n45fvjj9MC00KNB+uRtU8W7rBLuzlXyw7au70sGb
1K7EBkdsWHIBM8Ya3+469uRQxddiyAKb3JefUKnpAZR9SYlX/53LpCRxqnkelYO3s6AgEgurWAhr
uVs3FVyFgDKxD2en7vLSXvZTwjEjKSulUYDhUhgcOIkPFprRTrC/L83DvhubCu2gUnLDVHYBj43Z
qsr3/6DPh0EIMZRhaAfBblRRZXVAHnTcpRhxd2IJEyWceEupIZnZDDgrNhMYHPYn0yPXVGeiiV8a
Q2VMgEaIrUTRo/e2D6tKUFy9MzEU6jW57zCvQen/4ugMe9zML7hkRdFMY3eq389e4uRNg9mIJ0g+
+Cqy30KkKXzhNAUjb7Cz0Dy0v4A0QBKQYrS3xuJOBIKsr61AsurmlJfwIY615YzHReqc0Ba2YLI1
KsB8YkRMEt+o6ncm4jNjSJZr3CC6kHnlfW1ehDepXyREsbpTKgI4R5R+0nG6YuqiaMLYRBqkNd5f
AFDryw+2gEUBhQMlhlmKXgCOLc3VvbmTYEYHcJnxFgAN6CkC1c4Uef/XMc2n463MkIxjb1GYmx0u
ki4odp/2PE2GQ18tTIQWTK5ikV0J5rbdPA5FzxgGsqZJM3hQT//OVx8VRwdeRHHy0gG17VbZlRun
GCtftWqgpIa11kuHE2ADz+Mgdv84MDKk1n9ee70aOA7FD8+lrd4ww38bzUsRuPe/DRNo5FcXNiMO
AFw4fJkohX1G9rYLuFGrPY1M96IqnwWnLf9zpfTUCB3BM0YEhWzJ0nqdGZ48dAKNXa+vCrbi7m0/
qishY0m0DyJDzo2WkUvj5dEDaJainwZRdFJWPverGGJzBm4RMIv/7Yl5tE3LeZyFQrQhlhqohko3
SLJMqHCcS5xfvVS9PcEgJor9bEDRYJPSSsb72OS82c/LqKNRVHjd9WvueoaTSMl5u2vQab4ksMMq
DkMpzcj8Th/P0FXCAjkqEqSUf4twz+Vopgn/1+59V3iIxqEGzxgC0rzeCeITEvx84gKs6PEXAqBd
XvBU+eMM4z9sz8EWwlz7RwkCb5altOkAHC03kDqEUwvgPzy3K7evn6ISbSgL+mye2Sr78/ZtS7yq
sR3l91yGGp5dvZshbMr1j1PjHpZgNraR3mrhHU1y0WKU9MJE9AtskEVkYL5mR5k0Duw7vgjz+hN6
N8wSG1lyRxwbclzpK52Rlvd5JhhXwmhqa4hcdF2CAcAAY3O5daAHiLkBDFRZJ/5x7x+BprRIvO6V
a9yBfaK1Ole9GhE9psiD0rkjfFoS9dgpo0rStUTiOgAp0/RzG2n3QEYaTHR5xX51lL5prnqlQ0e4
xV6FVoDIkcePAMh+C7RYAJMJnsN01Xwi93S7n2BJr+7coDg/IK7zlHYpleHt8AS84SeIFFNj4DOF
kbdQ1an1g6ai88YleEuYXTwUGe49Tm8H01EDGhJzQpTPb1Gn5t5hYVl8Bdkjjn6rxyCwxZIPntCw
Up4hiddTvGu+emvjURrcLlmDWcfUNS+6tkJlH/CpafcVKT3kmxkNaIvd0lKxRDGpc8/SAHZigxpn
m1q6RU2aDuxC+3D//oIilfDYNVatB09GMrwbpk3ymM3eB1YyXm49sV8eeJUCq+KpPgJ3Mnp7W/BA
a6MHZNojJTdnQNalggQtu2NOOtoBbF1IT9TPKD/vDS5fm8fZj7ABuwaYgOeaZ1LKDWlmEEUey2TO
Kylv96NTPSxGoKfKo5x9iTfkgVr5Qq41LKoXQae3ECNWMFpKSZd7ydUBdJnmx0vLXlaX+hbZN0Ji
b1JWM/y90csNjNmr98WVsz1C20S6+2QQDbHNXO8I1BWfxzglgdrEv3bAtZ0e5PccvE3eQU4k2gVQ
2maJjv/0Tl4MNZ3rRL2FB2cSl5YpjLinGFrye9dxpc33CgAjNyuEUy7XiS2gOxZKYBAs+qyJihw8
j8WvQSuDJTAyKVuli/IBYsZGerIh7RBiZPRPKS7bYJecvkPshaUGxzbmnJVL8/MVRfffB91AKW00
+W+sQSfbbWWNlFKx1iGHgiTXX+Q8fQXR76clhoonQRU938X5IvTs36qd5hT0mxmsLBgppkjfHH8L
elcIihQeSEGglm7yXjbH0Q5F9jdj+vn4cVmQzVF17lfnET0HozS2+vxjxaJ708Aw4vguh4FN62HR
Ifsn4+vIEG54x6MYxiDK5aP1RiCV9YUCzqcAd9AOBAkTmenrOQHnnADqpp6TSv3SxAxMHPHU5kjJ
F95lqKS31rnQzoRy7iq4y/M4bigH0zxSnq0rfztezyCbPpazlKUKhQCg85Z4ZGpXc4BX0Cdxgcar
qVxyBUFjptxYdZ3h1E9pQympvP9+kr0MiMGrVdRMo2EB0v2jNosOwCRqZreAxpmXtcavKldxVBMC
zyP5Q0XF5NE1SVjhaD2B6cyfo4qrd0968ILuZpmSU7WtNWc0MOitYjsuo5eB1HgaglthawMWCx28
UMkQCcLM1vQBkxaDjN0jJA5iecj0l3pRB+240yC4DG5IicJ96hhzY4cLIUCxBHgnfj8lu6FlMIV2
6TV6lPMStCU8NpzOXSTFylk/iJ5LxfKaejNb/l0j0SA5SofOqcqFfbYsyyFGyf9ajWKwIooIH+/9
tMmdITQJ/eiMnBlu6EDDJhD0qff0bpfqoIZP0Tf9Uaa4ddV2htWuVZWtWMIcJ6fW/STWhJ3UFSqW
oBwAdKSjZEf+lBnJoJj5nyYfouQCct5/K0QAtYuZftvFtXR2gyoQULszA/g/OYhHCALtbFx5uUZi
DLjKfU9mA3aU149zT5FMzlfTiMtW0pu9I7/zB18TzGR6nVPYfLXFGxHgNQ1SkxHoKWgi7wGzkf0m
PYjsbEB/u2hIW6AJo039iFSKfVIY0g8iBt6QCQNfaPW2M4BJ4dEZzkU5hSTSAnA6lruRXrGmc6PO
1mAzeEx/XiGqcVuekvCq8Cz1H+2iTXeSmF9U03wTMqLZeP7GrgKnfyh7CLqT+ma5RnZ++Z6rkFa5
7vR5BdYAsSNtlms66e0ikt57Tdb+L+3zrzQJNKqOvb/+uzgYLpzBMRKcwwELJa4bULzK/iOAw2Q7
El0qiarmKK7dcHTDj7qSc+1StBajzjyHlBm7I5IJvdnI/6mNra77G2A32mV6/DjYcL5EB7qjyRLh
BkY30FgWm1Ks9AtqyJKbpA4wESn5LNZaeEV20nVlAH2TxbmqfaiT9rQYOF8eXy299gv8r1siuv8H
ULZ3P3/TtxkhKS0LXsWlvP5JtAPy8yxvmLZy20bJ8o3wDu/d7V+2zgF8w0/dVsxEWFfbWzXpZYFf
bpzDGtBYrwrlfiLNb1nsjTB51qtS9UCKZqaU48QKEEsInFsjllByBfnNsVskP5MER6RMEPxxEPfG
8n997GdeYfqFpuQjD0T4P1ZTKYO/Z9a+xuwsZyebX9q/WxmPTh2m50WbVZ3R9DvQMsJQWT5TnDzx
aQZgY9KLzMkx9Qnyypyi5jRDwMxpp4lIDSCWwdmh07hybhvczDtG8uXNW3mylL4/i8kxZ8elaxB0
fmVY+wj4I2rwp352z5qWN62IEx1K52kNXDgZhjLsT3JZGx2vQ6Im9UHPVhiNNwGLp7Qfd3IjbQQK
SAGd5BgBODDtiM1J3nfrseqkRCqywI86/ar8ynkAZMAssLMazEZV5g99nqYuUShkfmrsqRz5g5oA
9IgWjgPdqjphqjtlATWMivwccQjpOkzgaTaCmD8VA4zZLV8JZ2QOcX4eEyHmdQygmhkiys55Y4S8
scBQi34yjhk45YHwFbkxSxAseMzcoOtchq8BAzIA2/O4jRvrQdR/g4a3oPrDRM+hxFbL+9gfPU0C
lKGoA6Q3uqn92K2jwolhnhtHU+8/YCQ/MfGkhky3mlV7gN1hg+cKRWcUTbjdKS9VdCV0ijtumU5f
5iip5cWW7CwN3XSDyfXs/B3uZPG0Jzw85T8JOp+B7MKj0ZbAoDAjr+ozGq+uwQ0nZJNe+ucRja2U
qSQ3cvSzbtUyZNDs3Jt0tss36ZLAw2MKpRHuF0j60NMF1D7sBZLQiS7cxC+SFXJ5VBiHzPgOBuRI
Gz0JaXKWmrLipA3z4+Vw90PuLYtKAZM4h+O2A7N2wlzJJeTWd9RMQrqtJnAD60tigMOIEF5uXkyp
wTqU+Ohz6AZIeKgpkafzTszS26MuXLJTLsVJMgSJr5az4Gz1isFLmPsH8bDrx7pPKlkNY0DavnZ1
u7/1u+F4EeltwFX/Oc4znD6yhOE4Ul/aEQinRQvAKKtY9KeaV4T4Ja923r/oBFviGd+MIcIFwnMh
rpAJLDdqm5qQeJLp7NPV+MNxa9b4IPHLnGW/kXU/zWUBVERpe9SJJwWDndVNXfWILaRfcGZ4+fsG
3SIIOZZzBlMstIvf9H6SeFnTjNnqBRDHbnIgTT+iUAML4411GEEIGNfJD+YeEmkQPRnxZYgTCRYp
hvI39OX7RwyhmrgNdb54IZaUA2JBJAoJBWrQ4FUPGRIOrDxCATKZMUYOwGALfqTYONERnM/hCAnC
AOMjEZTbQiZxQSmbM5wWVcKHqvj6UTXoi6Vtkzz/rjRMkomLU9z+k9eejBquPtapwmbciM+dViiP
7U2HaHKnhvEOPIVkQ8erGN8OPJdUeOI7n+jx01RxdiN7rQ1A/U0KDmjRwndiz6oQiDFL5eaIVhjQ
dTOjX7ZInGa+CTgk0dtmf5fuo+KEbgNDBDAg6g8KjNTzRNDOCr4JSK7RMSoMBUksAXvX61uBMj3s
w0SXGAhj9+neGfKDiCipStgc1h0RVc5TlO3W1gXDQTjZcdupgGDkoXUxr5LPR/B5b45CuwIhLKfG
2AWrBTVekRL3GLWhYi9RLqPpNrFf4JnQKIeOpDQ82OhMhexj9rj7BrcdHGKH/oHGoR/onCfKunJE
/ohfgLwvdH06yURU4SInekN1XXD3EhJecvo9GOVmzlikGLTPVz6hIHIAfc5D1HILnjDkSdMLL984
RLi3VkyiM+7RA83jjZX58XyXZRsZysJ7DEt3wTwU/3WrAFJXahoCOw3/EqGVhjp8Y1Le8tEn5ZbR
DTp/H31Weyeke6DBBgDxfDwRJa4iZ2M4Y/GpR31A/nFRw4OsxikPe1Wf1TpbHl1nNgAyyxpmVUh9
uakJwasB6J822zskmwyJZaQ26mK1gA8+1Y8gRwV1EN1WesrLWC/JPfr7ZXNcbZh40PjoLbQZvrvH
lg9nDFbT25olg9kdXNOseQhZWP+D2vLOCwAdZUNbLyoHuLUctPzMxzcqTT9SBVO1Vt5SNcj3Dp/f
B01mK+eR9+9nhm+sN15lEC9a9x5I1+AvkHZVhnTJ56if8Hqk9ZxkTGctXfPYOOvi/1u+Y0qXHYUX
0ckI4A8KIhKzaliQkeI1ljl7JihmuW1ViEK+SidySrfmBnzs8VeCa7jni+PvE1LAxCXjJV9cFirD
QzS53sURqnDpilmATYyHSdy+INOjHPA/E3UUIvsUZ5Xg0EZVKpcbIQS7Mplsmh9P0DzOEDtR1CuZ
GthYGOYxnif5IBDl/QcSLS4nMilPhXiP74zQFlc2T2xTjo3QjCem4KS7pvn/Id7aajcFKpFohLkI
/lAKdL2IHpYGY6rdZaNRzM1Eu0psztm0Gr3Ppxo/r1gkvHo3CUI8k14YbCs/uvogWKs0lfkEs9iS
8Y30MJepAeOOfYCk9Frib3wKuMjmCZ8P59rtWkCIRUpDPg0YzXQ1hrkeYsSJssW907TjLcl2t96l
j3wEXqNqPCE0p/OYuzuD/kWgIzvIHn+vg4EI7seRSy4EqzNtTe++DdD3DBjDLzq9d+aGiIdz+m1y
QBKkf9XDKw0KTekG40bZ9qFHj0iEAn8WSIEJMbKhltrmw2k9zLXPxULdVoCv5WCDqCYaw8ovKBmn
qT1G+PMarldvcgAURHz1UTMKfn/WOQDsYBmz8KERjrbJvcKhOcibD/eWJaVyCoJqc37cLMKsbL7R
lQviHCaUdparZrsRzHV2HD+LMMoS6malE954r4sAN8FLXX19V85kE+YLJoT38EnttSpXCSqXPfDg
JWCd//gmx+lzL9rH3nw6t1n5a82GCXzrMmRCuYzfO+xzUVDkbrHD9+6Z/tl0jto+fXFemvcVJQ/m
f+tiaSutf+9Df4lbQ5nn0IsfAbu/H36SNia4IyXbTXoifIguGctgqn7hnJRiEA8qVfL3VF+KoYwU
LSsHiDjzBKQewmDkrp+fm5J2D9bwUx+avftka+M88SE7VYpktX4Vide4GRaGAF20E0nw2Wd3nAs7
ifTGwT6Wzcm1albodux7VVtY5Qw3BXNXP/hQRjZGsgO3hfYIIKk8twsLxyy5ejrhaTGEbjGA2vqh
ZjiCwzSG08tsUaCmHQ6RPyIOfmpfu7uIrqD9CIpXAjlQSdtd2HL9VDvdIyygXfiHLZufBadiBcMV
m0nt6IezAg0mVncw+rBA24jNFAgWQzU6f6dj6ZZ4Emdejr5yB3hxC/BwMVOJGq/tGJAkawcxZTN3
sss4oVWBG0NZ8tG3aOQoToXRBgmDYcceat7Hl2j8mlzwdOpod1LvU9KoM18kILmtejt0LouzyWG8
oAZEg6F1vNIUhp5Kj0g1FEKgZ2nspVyBKCqLYaIDrNxVzv2Nhpn6RMH77of/TPtWzf5BnfnFkneS
v/UgyJqq+tDw0iovSPv8KHjOLl8gfThGbyReOaZTlkU4YZdKc0UOUG5NnlN34JXqWnO0copsFB7o
gl0eOK5Ii58GuPRQ5iEU8iGqCTnJAbwcePwPjTAkAKQ8zPGOGNlXNNKq2m9eayDn2NWBvK5SeJvU
1IdAoawL0E+NMP+o5nMIpes3UQ+oWYlC/rL+La8bsS0rSW2W0Bb2vI5ot0t80s12HY9D2Wr1cA16
FCLaUxC0bsgY20vxGokkEaa3a1C2gOtRJ02017AIYkoWKCKHXzUX36U+G8XmERc+I+cSLPphveQa
/N9zMz2+38JCYMLjW6sH8t6nGswy6KEWPRFJ6NAHauEec39Urmr+NzM2OweUyFZnJPDnzfysMW2A
xTZPI6JfmZL+QioDH5x5Fj15nXN8qJHdjnzxeMoLfH6QQ58jre15Zm6bUyDiWDwmN+lrcoXCSrud
B4YB1UEun3A3SxDHGz7qvHyHoJcuiMtS7fpR9aP7gzJIQUnp7TucFFCeVTquT+HHkzoTuDzWjaAQ
EGId6JooJKa64/jmUT3+1MuLakC2x25kavnLmsL9+lNyiftfhYxEBWqDA+xd1hpnv8oZmHwvalmn
D45E4Rr6/MQAo+W8VjOGGssx9hseX+1TScqEfdEyEtYcxI5fUd52ZmrmgXHLWfV7NpkGGYp5biXo
x5B6MphG2xkNS0/QDVlIX8znWfwtjbw39jVI3e4G4kuc5Ey/9OwzUk8SWYRkk8BJTr0oivotx+MG
5Vo5sTSfua5SAp9YiSjSK7bapPmag3B/QzbO8MPZvt44XpsdNsBu0+vhIDqpaLnOF86TT0N5BdhN
REskfzXwYoozpcAUwE+201ApiA8Ul4Led7YuTdhrRaJyd55lP1D3K5XB/2G6ZP28aEEUVi0ZAEX1
K5Msoib/8+B581zSXGtxK206mUCHNoze2jMDh94RFDqsB+nX+qNN6OOA+VTZK6Clf3jYYPTh7JKl
pBgTDuDDuMsbnw37N12EscUMpz2CmFEctAV4x8KdhAIbtDNj3pUA8+G75v+ydhTfvW/TpP/pNi4E
KpyvwSoJ9LGiJBYNahJLOUnmVndp6BE3SFwPU44ZB0D3TYkIIPVo0iAukmuCaBEwvTE/guFwkunp
u8pd3NOdiMAQS5VTGHh7UhjmQswUduxyV/StSdGRbHZJsA/Mdr6M7wGWkQ0bdege0/t81bQ7pnkl
PIf9aOmWOoY6cCcRol5jrMnRgCGvv/4QR82/fZ/GvKoog4eC2NDxqsT3TKiFukB3lcr/tMBRqXpD
g0m9Vsjz514A5WRl3dXs/vm05qSMmOdAkLFdT159prP4JM09moSL5IN8RafkgLxHe9Ldk4gUdTnJ
T5K4r1yqzPDe7OcUXKbjs/R+BvrcrVgzZSid0buHQnrO2AVMWYq+93zLnT4Cn90MzvES+KgGRMWg
N2MgbiuG1CfqJVBhoBY7uOmTUHLgBwfbRvGbSn2zBidNjQTME3YI83AwU+NIga9Yykzn1KFM8MMl
t+gOc936sl+VjPu8tzjz3pewtwXcdUpLtFgYDFEnEbVCQkmpxbZLTu4jAumXaloJ4X2uceJbH9NL
aaD4ndzTbyVZxCHAZAQHgIxBXeO2ovqLG/xG+c+EbOmUZ34StrzUimg6LCybpuscX6k4KiAEf4f3
/izrjRi6/ypHmuNa4hc/a4poXn01JSIe0ArY2S9WW0qzHdWRw5e8dY8D0jm1G4qFHNh6/aGPpIno
m/vb+bFjk4jgJNVRdgB+xyo6ympcBiS0lGsC8rLlh1FjxLbUEw2waHS6fCwhgfRZmKDjj7NRMhvA
f6BTGoM6W5fM5Fq0tKvsSqkaKK56/TfgpgM5csIlM1MmcYMs/F0AhrgndziH+gC1hn6c7gEBtPk2
ZR/lIEEYRJVkDhbJQ5+lr7VuvxnNN269OQSlUvIlupMA3cI3VGn8zi9wRQ7qLpYfb2j5imCWf8DI
YID3SX5RizjQhxTFYC1pqelAurbAaJjcFxesdSOZjw0MeopxwXDbEIWAsCUgpBO/VUjO3CkgpLkf
8wmNRqC1batHr1SqBYTdHVOIeMQgLXattMNjurD8vByKumFdGUKZUK3Hx7JDDtkC0OZNSzoBllOS
6sC+k6/RgcQNzZ5j4v6XCBrTA0RP1/0gjUrrjXRukeVJDyBEyAhQDFNdnv1tOSH2oFJvRkdPhCYO
YsSZU2S018O3cEWwfjLkHlCP31NQOcVJ6bwN8KWti9B2TguemhtT/jSQir5e64w+iEQfsx14b6K5
0CeUmI4Fxh83C+4AyZIrtRfJwzN49nV2cRFuLSep7ia9u4m/IxuMqRKwDTPd+K4/rn+IdKrPgAJQ
34xWwZwPG4eo8NhWwfhn+/2+4b19Ea+PgYEQpY0ZYYweab6dLx212lDA70mKAp5dPTFBXSpfH2wj
Zi34IPUFsPOXTWTPvFBDVfNIo7FPoyXwNthHVIFGb8ZfmcxZWHNXOryd2oum5Mi/CE/Sqw0/FPub
LtRyxfYNzg/HAXoiJTOaqWpFWV7pqLXTxYC7EeHkTfHbBxgW/jWJsj3x9taIoUO53rXlwHLTupJ2
o5XQzVsdSup092lV3v4STrepQ40OX6weBkx8H6rMpyMPS9W7yjpje6Iu7P1FWB4MtS4ji7Xpg/Xp
WYr9SDsPN3QDSlePaMCmYzMm/OY1Law7SlwQghDZbIb5RgwdasMnM6txsVw2JT+ZzQsjP5GfH4OI
eb8cNfKcHSETfg2XKYETBweAWq/l85L1TXWgI/hYj7xInJjbXeqQlm3bVJjBP+p+eORSkGWgiPKQ
q/OECvWWwtguxsrNBsPlzjToAQowMiuNOC1jqwW3ASWpQAy6OJyjt9zFa8meGqjbL8MYeq3w5eHG
9ldakLMBosoCVT4g8jjV+doe50Ae/xIMCbQzyumbsf3kUDQyAVZgqGywUMaRQ5VEYlbEbl/PBh1u
EGn0qjx/T7eveEs7mI+vPn1pSKb7fejeZwoNao5WMrBDIKkr1ZA/sdsHlnrbW5swMzkO5r+qLlsv
tsq7UyeKt/n3xrq/KCpZ0c8c6LOfGbCp8gmYZFLD6llbTSZvJ371vi/SoIi2iUnFml0FralM3E4N
SCqHQfzOW+Al+UxZK9e8DkmR6ljo37F1a6Ut9RmlloZn/xR++A7jv1m38BiuCwuvW0CBDsTG9pSl
qnBAmMZXf74LXiVDCmFIiUpPGix+QjuI3lGmIZ//xniidYfz4pQnKxV/fGdPhmuzO5FKIPan2sqK
AGrX2Wzr/sdonXoAwKXYvGcLNevH8yFtFDqy0sopOW3ZWopiuCn/wlnUemhFbpgyNtCQqPANZZOl
ktQeSwUbkg7dL03YiOxUvc/YZZ44N3/oI01OaTZuxFLaCEPfVURP3G1Jcpv2qyoXKhBdaCqwGf/g
vIsfIwIB4+VMq9/R/8DqpW3qZe1PFbUId9VVZ921V4ocySAOTyStDEhm9koD56IM+ls5scVZTpor
JWRTUnYILw05J170WN+ZzDTpHD+jbUepZ/KA/2wh7YRDYH+qN5OCMEL9KGzvQ6/vxTousi4tq1+V
5jfjRnhvSN0j5uMm8e2H4k0Cfw6BQJZ/c/1/chTChmvXeljs04CucDXNW7BvY0ZwjEWOazdJzRpL
jak354SnxC+PCVoBWOQHg7Xl/zGGHhnsBCpYriQwS35kQXzCttZRGlrAg1hswbzslw22t9jKOWG4
l1hSUYOEko4Zx4tc05cF7sYlfyg9GjAw4a1kkOVaMbrcWgr3ox864z66bJgauUaYMVkdqORJo3WV
hDa/KHcIMMP3uaAj5+I8V9ciL8tEBuB+mivt9bdxeG/DDqRgFu4bpisLNNjHbch4hRT/m4y7MZrl
zOhHvkviABIHTsM/kgj8kWC2i7hPg3oLICrnOstObwwrnjdGCWY0tIHQAAuJF+tR6jxFC1pdNbTw
L8Dq7hc93/ci4jb9jvw/CZqkqWMVqPWBIRx9fq0NOMNKs01xGtEqufI/V9vIOgOYojY7Nk9TtbyG
V1egzGGQLVtzQL2nFoxTqJLA2IB0r0XEGxXcg3dBfofs2yBvXRcsRUONFJX40kG0rvsuKlYqysQb
pg+HzXaDYhQdbJerbnc8Px6u0msjq5Va5C2F/T0lyieAowmjZeRqVnb6W5D7A+Z3ILWEytbRjnKR
NkffMirtgNef8qTE2xGjfwePxysiLpEBYQdFGH80woAz7UlShZw3CNOHaQbTkKUHw9U9tkpVLjor
pxr61PMKNUTxhj/a44b1JX7p6QzRwx1DdhLCrh+Q95uJzG/cXyG2bZKdFkSRPP4WjS1LVPeSQ/ye
FsTKKrSMaFoyp/Hmzcxx3jEuH+HMOx53qRQRCMUtFLrtehA2N1kyawx6gNwD7daIIZ0zyAmwxc4m
i5fZb+HzGoHb2zMpn5DaXcIHB+axKVSZegX2IaQJxc6pU+iDW4grR5925DLm2fwgkG8UAyJtnRie
ghuCuwi/uDjpbG/UPlWCsdn0qq/AwDcyaVbbslzkyuNZcSvS7Kdtu65CEbaBpUS6I/dQ+tqz2KPC
CVHYsxvRcKJqJb6IRKf3z5efgwZIRaXaKYEuiTzGjvAUySNqDLcOpP9ygoZTTj3b/jQOtI/J1Iu2
TDilrMaWdMRAjG/GnosBS3HoUzpbCSBENIaUfP5+o5AzeY2JnWuDnVWrDvEiUaAAKldmI93Mrr9t
eOg6BLUVJWs/DHY4PoU1iB7HKrgTQFIj1ganY/UsjwWOFV+AB8yDHp9SV+1Lyb5ffeFI0dKP+qod
rlj6NseZDWdg8Kmz6FaabtLLu2wjBxsEshPvWe+KkSfv5frt1xS1lx8zhtMizubgmSoj2iM2Qy2s
Ee1IYSzSLzB9vEnU5fgQF+QmP5ke5Z2y+SeRkN8z8iqJbfv53dxEPuEGyzCVATDfH9fFa+lgyEx4
xP2VZqiNTyuc3/asQOuZG6HXSZDfkPUDU2kO1HryKv9Ars9ySfmqt1G3VFk+lCfWt8AMsj/IKAh8
Ue3imMkoWqPbsjNl4kjiT07YjV9iLV1ARyPCjU//Va0bBY9f/idne/0LMycjIuFReIFKbvFkdamh
UHR4MseexBS9u9XMMlFidoaR0J+AgyxbcYaiNvpCPUOskKEHj5sa+AmqKeN8JmBorX2jj1hFWoWT
asNpRTQjjzmweRybGO0Uf18rZcg3ZV3HaK0gFf59ycC9W9jKT9vF4INq8ES9s+VTWiebTrdtSBp2
IMYdml02zmlICH80rwZ/+bmxr8yITapG6soKYwMcAqfpZHN6LPT0lqDXR0pWR/QbeYQDYGj7J03C
nrHQLi1tDxcqicD8AX6kTjkrcEbwO+wohHFFMOdrp3gbLXUfH9IkfIUZKOoKgE0owG/OdRUCYNr+
8z0xD4IaOMeZqgXnE/mJbFt6IUjhLa+jbOK+Vl8TXmPvc4JP4HXr+5hmvK+fZYQv8e3ZLYUPVCbL
496QgPgK3M1mt4RzuQqP8V+W0tqwDJ/wWw9IhC10PWau55f41UcwesQs5+3FN2TwSgCnP6SBN6QK
+ism+xaDqaUTQGkpmDsBzAeLO2+55nw1Jiov48BqFlmIbwWUYpL8ZJ5ThFZpLn8Hhn4A4nPnku0R
I9CHmeroxd9PDCLHZWy74g2+Socj6L12K7Cgs0KmkUH1SJ+S+8SWrtKyONWd8XT2YlakJKwUz3oU
VXitz9mwuC+jnlGjVEXaN/ffZ1dlrGsta7Sp0OviCf9Iy2etfgVqxvBrxEDn7o7t0n4UdZFshNVP
pLMq3CiIBhsl1LYdxYgBrxwOgrDPoaGeXKsouklHm1nkRrzdDy96VUGHTZgNTVrY4pLksC/a0K16
tqEu77WJqtDfAcOEjAB98icSa/2MzMihc9ecgkIn8+nU4VNIjTWs4Q2zJlqb0dcV4izrd60B4hb4
bZlNkU0I+8UUOiwx7P1ReZyNMsL10y5gOtB9HemSW23SUOKR+GT23ZwjZbiuZ1C+k88RHw39w0Ca
VmGmNa+crK2JNsHYgY2oW3rDc7hpCHDo5aUpkzrmjd+aM2Pr4YBZQpmj06FomB3MCgIHkIwIuJgc
4l8rpnLDVDJUaN66JQTrTFpfKvK540DRLAFP9C7/3Y+IqrdK3TRcMKCkbIyb/eQbq+XDUiWwDlj8
zqs9hvVBK229YnSoEU2wweE9c/87mBpxXDOBQG6kp8qLIAqaK9z6lXyBAifYfZGHWjTEGFeor1r+
rm7pEbC1drwHleeBnRciKltOG8SJWAx3MdZA6fx5tTswNERPWWnTooY5T+qNS4/spAvLNC/98Be3
TRTpvOhf3wpveQF62XQEz8Bu/6Vw/A93HEPBk1X0lBnSYztuNLgc1aXL2NT8fJ2sltJn6Rz6I8Uh
TCFslPpyjEdSRgMW4mpt+f8odcUWP+j26BPWl6RExs27ZyhDUZxM8nt/BMC/6e1DGnzoWCNvxv3p
nfM0nFERugEFU0OfgiNuJVtO6pEVubroKCvVKBSWo8sw3307zJSJG7akG0Q5xCwPpytOAmTVCVEC
IVSoaj9c5bc0IGIlPtPBgzXu6e60rTapI3hFUuZEHt5NocnmS2O3vprs6xjFtzyaWFh6QFyNRg1d
edF/7BOBTB8185JELkBzSnlUe+qRqYGKEFV4/zPC0pSIOST0J2a4212Y2UjFtroAPC49YnPem6XR
vtjL8OApzhPbKMTzjmuMxtkQTi68XWcqnNmJFyhVPnPYUJ9i8JnZbTQZPxhsxL//vqCvvQXG4TRv
OH5zAvEvOblM6+pF2Hft3n/WFCcIBDnHwwv9TirNzQAWG5gKnV9+i0DqiTl5F43hgy6KE6EbwQVw
wdys97D7+5ceRl2tqJYfNKZKKJBHPKQXAnfQU42gcWycw/lo570temIOM2qBJKLx4H1Sp8oVf2dq
AE32xIvEPMxjxWdANfqd9WlvLW0hoQPZ1vQc0oEy+MiwkPfjIuQe+pIelNsODlms2e9B0GB+zQ/i
3RcJZ2yrVAS2K6z/M9OIa+SN80aI77b2B+8F8zWW9cTIU+Grob65RBBAiew4CyUBbNi0Nz2gIlGr
2N0uyIHorkuRXGVmBEiN1OhFKgSiF9yaaFGbS+KuAiDt5qUJoB8Uf9f5sU09R7R61TVw/lUefFLZ
bECKHUUmGrRc4IrUMAEkpq3CZMfFbjHGJo+jb0Zz8EmieIM5B4XqKLxsqvIjamwM07pzPpgrFZ9V
oogazRVdIf4SYEawjo89Q4cTFAvx0oCyT+ky0LOl4fyB6D7TWvMM3XlfN6ywah9FrOgc/BZdsdIj
Qc3Tmppp+UNs7OJQj2m2qCRE5Ew+os0TOnS1VSz3CpUibYMwAHXe3eclaEUdR4PnlKps4KIwa+RZ
bEHLY30uQe7p4N2nZmxU6z+4cK99bYWQXJ58a+g/TVPt//mQaLAtSz/qCh0KIYOqHugajHhAnlti
SITjcP1rTZ7e8r3BMbVBC+3g5tbPSm9bh3cnsov1O2ioh+P/6f9tCVD19kCAZsAXJ3SJ9vmVer5a
E8/t8YX4LUsXH57qBAypZZXfckazO3dt1Cz8G7UiZ9LqoAzlHp8XCBxNOjuBBH8NM0RsuUpFJWCA
9pwXEIgoPsp6njkNKw0/WzVT96DLJjrcjOa/4EfR5KYgBl1WBV9oVMcVflRplQj4i+JYzoXD8Du6
MirV6chcKBYITTFYSEhs9ay5cf/migsVl1DvZ6HHfRkDzWk3RKls/76AZrzqR8Sldwe41byMWO8/
g8qryHIqkeFJropZSRXKGj1ZQeIXl113SyDBsDRrdNeBvy67M0iUqE9KzmQPnSeaYgtxoMtVCDNT
HVs92VgYEda4rKjOKHyE6c8hzl1oLT+btUv8MejSuIY4Ojy4XnJekpCPowGcduCHE2NXSq36v01n
wcxoCnQM5q4HwJ6rPuClAp2veqCDp/cL+kkEmGly3/hVGI7XMkqGEry7eoGLZafHA7rPKNVPEifu
Z3r5Z0xoz/uRwP8ObFK3pgWINdgFhv6/0bZ8NlUrUNvLcAqsmA7ct0puiTTMSdgILY1pQcNqguHL
a1qUn/hhM+lxIYuhizXclXbVGnaTWBoXkZWpGGkdvRqHGlZT85pPszugb2GFrPugXPVSekCz/YO/
8RUP27Adz3S209hQKHbEGJey/HAyZqCB/MkChrD7id78JAzcCiApiXMIPrmCMBZ3rJTnBA8ekg+v
7RmEAyaOnIn80zj/TDfU+RrQ6HeMNswE6tcIQBmMuzWbjz7p0A6/XBfniVmdw8qplHr4WEkyRwiH
gzqDpgUz9NkQDaygNcBTrsZIho85y+SMj4Y7kOl/3Tmct587POLAlj+Myy0nn5fKhS3EW1/CnUnU
7jcocbrpSR5JLnkNgiafBFFf7SvvdT9sI7Ysa1DNWqZjgQXbtCa/XQWnLlpiqjz3n15McytKBlO9
2LvMh3RXroLf3L4B9K+8Ny5hdG+qc39DnOxviD1Rw1dyQg6Y/J80E9aWrUhLhSWZN81cVWbFKW0o
E0tJjhX8aMUx29RARiMbtgDuZs/rJ6WNBL1o2pUdK3P7C+vZka12QLAXU68OST5oHgjn1t3KyK1M
RjMABxSCTbVxDjD1a0h2VaAfqY3hIBmyEN2kJyt8FjVguRLUUAV8InUmlakA3dRpZgEvQXss7gE8
86fnIkKW53FSm7Gfy+ofu2BU+am8VCY9U+EbYwoCONrX2m8AwPDyoP96iwwZNiZsCPaoFeV1Ty7G
h1aBJzKnFfkCX+pPMqnYP5coRCjss1vp4ifPQfmTfFBhd+/ZfWh3gkzfeEFJ+jCB5Lk0qrVYBHXp
VcjpoK2ewdK+TWQ4qxJrHVgYC4OOb06FqxQeqxBVVB1koFYm9XX6Yi4As1SVpbYgdN2HCjX1o0TI
mi2l8TT1tYzeDAV6GxnLSWE3UWfAe1/Ma3bcG7+Sasld27JSQzR9VjPS2lCIedhwpvL5g8OSv6Y7
b6IxiRuSjfhKIu4t9B7gKmgrFC1S3X/dkepWrrfeMawtjSOd31Bq9o702zWE02P1mlbugRQ5mFoi
YqgE8x6vsORqV80jXd1rAVN8A6J+aVY7ZMbf6WDy6ytVm+yqTweFQ/Tt+1a7zZpxNKiZ1f/KkZ0Z
mlEjEEkD+GvTnJG27fE1K++HI9gzUwsV2pouyP5mXQeUQmKbG0qz7VRHOd5M4gpP0f6/DNC701wt
cyVjWdySgWK35FfhZsMMf4THO+G9KQreLdJqFV+bQ/43T28Fp2bfYYQs5hOk04STBOspI1kcCeZ+
0gvfEVOWMmQbpJbKlI3y3GXT/qi93cTijHfBClU7agQM1SYQWwzRIHgQHlNCFUBlGx62Xsxc5TMC
lEeyH7jHgh9yRTTDjRSzImOpIVsTOikqmdMo7E3nwWXbT2uJiKlSJb2cLNvBRQ+SlYBwgJIvYzRP
wFilQafOBlQujFR7N4Lvr/eKImnNPNkKLkytKQWmXFq8OL5pHOXLQHOQykhbHm5Cml9B6OaybLCR
rAeAI8khgqwYNi+0FRmGUoq12Ursp2BZemgPht1bRkzIipdGYNvHa7NFR5FvVVHckO5pPTb6Up81
uMOc+ed/t3y1pZ3em9XhhN+u3pQzYYwh2pAvh3z8l0Ys5oiZZpDSfOgVP6Wwm8Gb6cPxM4OD33Nk
g9N41UG8g/gIhJRl65f9FSsqejZC8kRlTEBcVPgxgXUhKH+uWCF949FdSMFtBqDNFheMY2MDSihE
BN14uFHizfqaU1fpCDA2KokKwSIV2oITYuLDsKqXdnaoj3j+hr5e/A91Xp4jZ5e0j44frw8Rff5o
QMvOMJzN59NofNkU/jrW62OQDjL5w+cdacpD8adSPImw15zQ2TGCbMiYAsVA0gau3PuB8ZY2KuLp
ID+0Q8sYdxyr6okVgumnskjnX9pbxkPt4j7DFr+Ad4RM35YUlMBubZdIFRMGQtbfLeaTuDhguVyv
OVliin7AdyRtN+NLFG4NVMfP9QYlQ2BURVRJ7M+kQyLAtzdJHC510vLBhN3dFB9vUnFJP+sktxQ2
NCmr/BWvlY1fN4iX6nYk6E0zZoyHnsx/UoT2zxO5bHkWxCpNCSr3i6wFYum+AedPuOLvvJk7uyrb
K0NxB6KpWFfe8jGiLSnzzI1DwwjZL1UJHPIHhaQNcScoGpin9LUZr41+osq8WF5CNtw2UueZXNis
rNxkOducP7wpJN50ei9GbnrLH1rvkfJjfIi5CMMVvWzveCqj8DeXasMJnVd4PDgw6n8wrCDZrLII
U7lfyXKz+EojPrh/7yGqzIvKEh2ux4j7Nt5yr5kiWvfLYOJ2N1ZVyzMp0SJANk/pG1Mj+/GRx18L
EwlYu93JILypFLrljZ6YeKfzBxWylPDWxKhvQdvBBa8p+bFCM4QBOB79XP+RCRlwIQFybKk920wy
U4MXmJgOfL+v21cB2JUqI+fyGLntq6tVWIM/q1LlLA9I/bjYgW2SD+6H4Kaw67VOt33WTnjUJac6
JDX+DI9FdLm/JyIvnMDcbSomn4jsSjxNPASvpPDhzgO507E2pnSjiBI/bROsr0LUMufchIO/HuIi
Dtt56kljFdgQ09kmbP5lWqIrR+UN2JI0Tt+jDPGD/pnKzqd7B1p0fHj7lHBlN1FEiZpYIj5ZFyGZ
CNANTbZrudXoA7YNA52H4e2w2nzWjSzJ1ecrCoFySyPYDWi4tYfkTuBdVtKgNwiVhPCXa4S6XKxM
CBAmfXP52k18Iv3VIxE2LPF4zpRMqy+QFcWEpHJJmDqwTSOedYE4MYkHe1FG+onYr6i08R9upZ14
mh6xUWsmNMZM3vMGHQvIn2xSqO9hTjFBtSMUjhzGixs/YtEHY7CPamuTYqqTedAg1RVOvT4WoyYi
4pK7/Cj4rvvIVixmsuBrARHAQ1jg2jfyrNjpNZgrW1j24UxvMSIWyxGg5bZpE07+IR8wf2Avjd4J
ADp89QMbdEuSxglxsxIDOcsosEDcIjcD5YdWlVOtBwPhaRLihbflHk4FP4E9V3XYsuBljlo3PERa
nH+yx8KKDLbW6xTdCRXTc0hYUB+A09OWgUOjkVIEUtrBVrsU3AxeMeA4g6vZJotCnVrD1dssjBdj
NfxTdK9mwWHZAtj4N9KAN+sp2r0nZ+alIWfaAFBziX/a81v99hAIsfhs+DXd/24c6hCPall72WGB
7L5O6i+NevFKOmOuIU7mIeNxGL0hFnuDjrlWH79VMmTb3GOiR/bpXIefYajuVbn1gAtdq4gNzbcc
aXWDeFl6pWKpu9MrSyEgJPZuw2BpqRHU/tqCFoA6RGfwqZd5DUHa59P5Zy6HW4CoFo1zNEn57+25
j20HBGS1yKwWy5Nk/93AL99CEQiclpzrQzOcpZT2nQuTJwEuSwIdyEixkqXBX5qguVTt/5sfIryq
tJAx4BAojLdjfvxHeRf1Z8uPSCvq/O0z4AFmvPgvfCZDwPYctBwjpG4dlccBrpkz1+s6Gn78bLOc
VGjU9KDFOr2FXE8Mzs6mAt381AiHQb+25bw0B0WCvLljZ0cVTipbHvUhf+W6sThFJK3TSLmXTmcU
PHL5NawXYS99Fq+LjteGoqPtZM/OI8Xu7kTYxaYUEhiph3RxCooLbYtowcTM7LHEVMeNyyjEnJZK
JSEHPl3Y8ItbZPCa5HjPEzrswojOBXQjFS1fNzaY65EATkcYAHDJblAHDt3Gmau+r922LzwhTPmu
5kRs3lnko4MWxym/8aZUy85auj/drObvhpDCetyV9/xFFPaIwQlcTnm+M7dM6yZZHXHR8OBfpti2
v4hhVFjZIwZqDaDXbS6pSRXdBfqptwg8+gL/g1EU4qFAZJNhgDn43xFRkOqaG3DMGvkJ8ThPVO5h
+GlHy2hk09Yu5ZgjwFlEO1fEmATV9EXwn18qMnpUeJ9uRjzkt8nzjz14FqvzfHzoduJ3Tv1OhjVg
VAJMzkOL6N66o7/HCLsxYvtwIuFSEXKyMhw3iy/4KVdyvU/CaJ0fkTs+y3D+VEdU04XT9MSfFA3U
/5VyD0ejFYGb7SpVnS9tnd5qjrCNFJPBwPpXIRnxO/cVM5VoobL4DBSP4kxr/YEGMPQ3Ou/rJQ7D
rT2l7ROgkKiRFQQv9utL1XlX7+TMhxfWiTcNNKo8nR3CXhYQ1p8hzg9YXlRm95DHJA5hNqf/dSbO
cFugqHNz8uL4E7dOA9SCtKN7ShXwnUG8BRbvr7NfxhhAXmE3aTXX3JOUYnRy3d1RXDpxbnvlbsuP
1zX6C36DnK4Fqg4yzojZHbfEQHKcNN6xYvG/vwP90g96s8fZNUOmNv0sjwVFguumlJJOMu2Oqvpf
KyAMJxACvlJ3MuGYPMPYMVgXV1IOtOmVk8GDMWUXXDwcF7wFuKpo8A60bXrB+8hE9T6Cwm1m3ezD
9iAtOYmk1fvzSsV8CuOrHl3siZy2GAKd0zbkMMoTQlJwYuNegDYvdZWThYKy8viWl6JJ0tRzVzRu
Pa+FZ5pJXnFjNvd1H5VCf946bwLwCVY45PShBAOskR2JUy6JXHKp+wQnpaENWQGmfExnPJQG5v7v
di3NknlQWSS0Uv1W1peUvIdbPmgTM1VR7onVqxLLABM2TuNxCzQhHsqvU28pOJz9Wd3B/GmMTgaI
iiLTdV6T6/e/9umkuYOlijFk1b8dk3R4hl9+FvyyoDsaRAiBjjJStll4tVFRRL0pcLTqzW3Fw7PO
ZDSqFLHZ7MvBfnFzyvdZNs7KN4bqXcG00d405wWQfv+xAmJizs0h0qTXgYfkw1U+1/OKLoHXRTnL
Lekc0PqXG++5Uz+h6c1+YCZk4yNmwvJH3Ih7cxcUrngLw8ctn40CID+1axW32L84S7Uz/+fSsHQn
PGRhtcvyIHV4iAvO83xNBjSsSLv/tyKUS3BRBi7yigY3c46Y4CX6O5eVMfJGYVtFpTuaN7GDwWff
o0DGsTIfQIxWBFklckiatKvj1K4w/3HeuRTa9HR0sTDxTu/+biUY50QoeLhVqXXdB7NhEQdhB9Vj
imSa9iISGaCG3ffBlpWiO5f3n1xbibRA5OSMhrJ1oAhlzt2ScNqIkx1bZ2r9th6sumC7ZKU92eEU
e1r/vVy+u3ZReSZQp6sTVN3H/+YedHxxlEyrS+yHxjsdsB6Tkgd2UoHS49le7QB36BILXkgigzN3
7kOPe3RAWQtHweoLxPzE+T5RuD213O+edVbqQe4hN15tgmISRH+QAXWksith7N5TKzpeZo3CMT6p
xl2tv2vHQGq+O1qkCyhpKdEMIgWvGzLtNxP5zYwFD3oMRYBWzr7ORsWxl1EA4fHxv12qP8TfIc3M
9SPu49OxNH5Agq7XFGs4GW8gchcXc0XXUNvAvMxx3gowZwgskYbHntirRwZzldKRW5xliJp5Dq1N
twxS2hF337IMztJLM3iHS0MTWM6bO2vkF+CHdht9m1F1FmpmrWHXQd6eXaMxXFv4zm7GvtGYwxce
TTbxa9LXYzb2dI5qGRw1Byra4hfdcFSXsu6PsGaY/18oTiiTYIh06Q0digwxV7vKIWR0DQUv1/2P
wDWZs7lXds03gXq+Xq6ORqu4oxkWjwiMdefnV51VBdTFvpMuwBfDVfsY7ulnHXX8p8TD6G3MEqlL
QvzSPMbmzC0QsAC4cl0aj3i1r/fYImLxmy9X12EfICyWekcXmCnAhNo0yfVnEdRB7v7Cspi2AJ0l
57F1tWsC2KFECaA/jO1vceNmFtV5qanFCBnJ1mmx5Hd9m4xpOHhUowQZoQ726zm8fUNPJbDdhGil
IyEV87rpYBehOeSai9qIHG6Lzsqrz0t2f/Ly6t7nU/7XkoJou+8Xopf+IaKV7zsiThCSrXa8Njbm
2rDtYPk7Lj69CmSTBkND5VSokNbDcNldeI6mwXfhbQi6Ki04McJBf50XUQWEHtBFz4URLXw978ZC
hpy/q5FyGJie5VSqW9dcpOKg1NiEg9Nb3omaWC6KSD0PVSHeQGWpfaIHNosXxz38d647O2HxAX12
IelB1mJ+5CwlXSFxXFzoNe5VppQGJ8g+aLwlEK53cvNhvxTtkm1MF5x5HfM3VigDf9Id+pchJNdP
oywKEpqcON9rrRYAoWX9tiDYffNpfbmmFokQHHdfY7E1S9flgzz5S7OvsWkYUbLL2oDl0ScjriP/
HRegu2zUFZXxdkZz+PEcbisgzQnKBwUMYrxEZY9MApAGa5oJm1slgP4BQ7xY/G7fTzCtmWu9tUsF
47IAyGzRZRX48kpf2RfPwM4qCH/0haPRCtCm3RU3u4KmzmoidX6U8pvc7e6JDaSGVnSzzgdZxnZn
DE3ozry7fy7GCSXS7UyNTHNkT4/2TIZwK3auS1G3K8XUnKe8fa5x9QnyxXQB7r7LG9RgP5kCEkpb
ENwvY51TxQQhsX4SMLzhETHeKGbNovkXyYpXG3G/ioiO4UUmCoO/0SubG0n0cPNmXpr03imhmP5d
0+blL/O5H4g6ZRTWdJxOE9WJJPJUnXdqV/OmcgcgnIOMsd6MXMmGRcikD/F/l3YNIVb0mdadS9FA
hEKOwH/cn7XTshdKbJUj3T1AuIhmtAHIrRbd13XRdVL7CjQtQw1ys+qjY8vkBDhcSNDongixlm9f
oNczAIodtCLuY/elunDoCePly8XY5TMUwBTeAa1Qozz6NPe/5mMsXaIiW55w2NDun87q1+iKdRET
/0bq+Ba3EDdzSvxarZ7lU50pUsVaJhwkVg/e3ZFGK/gaxpYk2nVGPO+7tlXzavunkOJAk9c74BYp
Mdo2Vpw13ox7dzrgtu5gvhJHH5dvDNqANvqY/L3wKv4MHkMr6h//GM9RbRTIrDpQxCECrH2bE6du
+PFEJRlf6Rzo86kGraqPFFwM7rw0/6jMToaK/tvJOsasvnWqQpebSEEaZcMtyI3ijaZ8eK2BIBmy
QEJAdcsW7Q5iUuc0xz7FZVYM4EFhvlqtBp38JcKi6SB5p57lkPew/D+yewDMczOuyvK+uigWbT0Q
vPHxu4ISy/R5hr1y6RDeQYCu8yYDcRw8xdHlfDKVDvJAdutTg19YesymotKRicp5pMaUL1OEtLMk
9kTV/gkqPJP6apTzqNi3zd56XgvPLBPmMYIOOq04OqNCVy+VIGIIPVF7M0gLR2NkbM0z98AvyCSJ
YzyKvVfHKiz4RxfROQNWvccFAdjEENk6GTa7Euj5cG/RliPFp4iZLwlJGiSvb02UsbBtIbO4Jjii
YM0Cf4pPBeBR6NaOIXfdWGdtmigwAjVVnorrVjBeida1oZrbEuf2fHO979gW4k/bVy9UuX+jYgwr
N+ZWuBht988c5BLGxHt1/G4fCOUYHD1c6EPr1/MuJBaJTDyTFbkDpPb1/60IrSuTdFM/h8192OSk
y7GXt9+CxBj/RtPpTzymD4dO6z0y6/6LFnsQsCsl2ijZ21vpXAmk/3hfDaZ4r17ST5rkmOSZEg8S
/Bq/vHCnnST9g7CBGjjuQMNFInNcEs4q2QelRPRyAv4RyxhJ2i772FsQZ+LnQyUiNWarQzjxpsd7
RYZnat0wzDBX9R7bocIjvMLYZuurPTF8AWf08IynXh/oQ5cERsrAWBvTVigCUCN2lS3lWYC3XmjX
Fhveo2OdYFOaQOJPMsuYBNbg9BvqNM2T2cwaznsvyhD3xWTYRmqmxFnxcjBvCzKpaiEJZ60mohc4
kjzeoTBVMTaio+0Plpms8ADixVSChAjk2UxNxzjVNL/y6eBugCe26UjVPjUGKHCv+gSEJoIarAy1
RzPHdIzg+Y2brlI11IC/dMoEiL+nJpmLvXYbRzMhOFi34VN17SkTK63VcdI0GkUvoxcda9aE2b1Y
5trM01wcNyJRzaS6AXrErVIn2ZPoGGDuC11RpL01ih0YBqsdzb2IPmtgQ8AvtqUc4CV2ajeWYHk7
eHA5fntP7LcU3DwNMxL8DiW3CEzSxxgfdQsRxbruRwklBl3p8hHgsrx6JOKyWL0r+ombR1hHjgrO
Xj8Zrq9hvfhiE9HmldvaCFf0l06qeN/56/5xsIhK7FM+bVAUf83GwVbWHLYvdVshBaYPqqmDx00h
FsTyemBEb6zlIZHfkeRThXWrRwh2V9A2TxhtQpEGDxolsjoXgdiXR91RbRpCr10H2TKrihL9z4jf
8rVDiyGQx4rXAbqO7bEehbb56bu46+y6XP2c8mE10oiSiFvdLHiJyC1pij83B1pTTceBaf24AIc+
dtmPNK3JIZXhcz1SJRq0Bcc+SRyQh8sL2xELrtg+P9W0IIyMeb1C2fLLzF2tlLmKr4jWH4MjK1v9
eE+ZmVpmqFK9g4kn0rmqTZQwvldS+6PFCKwgi3KQm/3we+v7FdrC+qOdtjYEL0r2PMDGFTMTxAWC
SPmcJrmv8OIjm5Uo/J1QneNVeXM/evPZRfAkcM+vg30RS79pWE/nrcGCD4s3vyMmmK2DOdqTdBtX
hOuGqRL1oeM45oIexA4bZdFKWA+FvH0ivdSa1lNRzrg+gzrmudbfRoxLFTRNrTQzL7EhuZ4QRiYW
0SKuD3+0vW+8DQYx/gVkqRB+n3GeVoYe97hDmrx/xsbjWO2tDiQeJtUURK/wOGNW7Bi9/CR+cNKd
7SRE4EP+h2z9gs01yAS25yrTCFkSmZEv17P8RXZFJHJV72JVN3ep0JYLP6nc/R9cH8iSmUnSqN0D
0v0/VOEI/Z4Avt5fg3CZp77Byx1FOEOUTUv/4SxFJrH/Kq0cKChr77aYRFSTLx3P1hQBX/BSwxej
zjd2o36fdAUoZNWlCrkriJPodh9ZmqtUrb1gSegZAXKSTViSX/DSVopkMCwPgHpjCgQwYjBIAGCt
fmkibouWmlB+iXamrStlkqN8tOas7E4X58NU0BwIpmL6AgltAfzqLCdmSIJpiSGNN1eV/G6wQ8ro
qWoBMeG03GDmPKfZ15pEtCpqZT+X1PlaC/8S/ZnToZ+iSUvyXTcc1KVHtKXYGmBknvWb4iH0mjKm
WwiLdOCqxV6I/QI1ntVa3GjYns9McYINIDSAd0kMgBmGceRAVX1tyeCOpAQZm0ONcR4fQkB/kvJF
IPlpC8tHiyeWyT4ryvC65OQhjJIBAczlhRdacd6AQsRvQjq/R4lR+6WTb6wZmegpxp4sEMczo4Il
3Xw6CfZ+JPPXdJdIjXlkjSv9F70zG+7dEaWr2yigMa4KMg/vclpjNwlidgU0347PnhbnOEETFs4B
KT8dgtpU/M0spEv7D7tePp4zy0b4/FJCQrFfOMm6tc4i1jCcXA+Z7Yq4Mk6RGYrmz/2AUB4pzmts
Lpl9bqo6rpBTIFafFiPEm206L9ZJZPjHGsPS/XSiUlXafXkjCC0NvMHDrKCo25PTrWuWJ38LTRbY
Y+X0CXmScukdxsa6NbicJCg0re8RTsnQefjg9KgJfWoFXIDN14DPyKqJHM3G3cVCPdF2aNsvcTCd
HBZ9ybTxRzfb/ADRSdg3eXqy563/iygr7fr9fqVnv5Ke+pahUNgwN7xrOKs+T0X4mwaw7ILlGK96
d10pWP+cgO9yVxY4FsGX66weGOAk/yIOoU5s3gfOUXF9NqZuzqzp6FmkCPJSC63MAagklB+ft6kp
Cn9VRIQTPdHIpK8ONhskVBxCKRz4BxhcwpylYk5aicFf1r9kpXC9EVi2tineVvuhauXCdzPD2OFy
sUZojt7BN7ErbixdxPl55WbDpzF9wd4dEo7wY0Mj1AGuN19YKL5o+aer7cPH8Q4LlIDFsxnGtciI
CKbg2ddTe4AYbHCK52L3NDOE/XpkAaP6sdXU3wSWzo8ln/x3mr/d036s6Doahlgfus/SpTupeCDY
ydloyRy/YnRqnlaXMG5tNwAsCG3vVIKosF4qjOefrxjTwZrKc5Mx7Brf8d6ftZ82KFv0/WFMm2At
dDyiRHsrPSLoHgoKCnGkd1M4+XqGuJYkKHrKcJEljWqjXRbR2HoJPKTC/vdd6pRL/KcsD2mMT7Au
QFBFcVcFSgzYf/GYjbOD/Up9I7VA6juFesO5KBqh1LymEAKxAESQ8Nf8ZGPKQZW8GUT6FtgZfLn8
QdlOTefYhMdbSgI0BY5OhSW7/0JllnR15oEZ9bv8AxZd8Hlj9Pyi4mP4t7fvuZKCUwoYcg6BW4Fe
CXNdIPQezGqR2W1J8UXmGBzfWO/hGEG8qPVsgAeFvp8tvh68yPtjl4DPIFSycrjs4ffICZrJSB3W
NfuVxunQPLB+cBbG131ySFGF1Mq21kUHuedf7OBl1azdtYEypIDF6GnMOK9+bam8eWoxLyi3ssBY
5ff5pQZDuvDYBcU7aqtwDFJabSL+l4IrpNMt29OsJIYUxAqcro0dNkc878j3Z0K+onRHzZRnDYbq
6+mHLwppdLvhpPkRSzbAx9Mg2VWjfHYTr72kl9NloesY3zxGUIb00p6QPg71iHoK14KyOrINFqji
Gv9i88iNRza6aWllEaTEyE6+hmU3w3UGS/plPxpixMIexYkDO6ge13Iefd1Pac4AxkoX61l/Xj0u
EmAW3deXFjr5fjxgXVNJC9Zbpo/LHPwxIcVc2CcnYkAdG6iWbnireffLzXRBZU5Z/gMaY46q2T7l
6CQ3t7abtuihWdaqX7kEMM/tHfniSyCYT5bPD6xXbRL5XG68eIo3Yk3OBDR07Q4I0cO8UMxSgMFQ
RJfqAE1uy+xIsNVXy3HDpLm5BNkJJW+cpWQP3ekKefWTzjSY3KKzbe9QwIylYBehfc5pTBt7ErGS
KVWrbcGcNgn2mU7nbb9aBuAbSSBr+sSnRPUGpGx5kleP511CHavckr7Los7NdbxJ8spjeQZSixIb
X30fvngbETttvxqQhE5y+HsefrhwDFuC4sy1KtdzAEfsqLvtHNU6IlwR2x+zIRdzoQrwe2olthSe
3DzzyjVErolLq6Iu8gQkr6SCZ7Hn1Ob/n8Dsdt8HPJv1GnRJH6y3rsK6D0lx3IlieDUakV9qvz/E
jTrnx00hLVPNlr/x4QG1SO8MWHF6eRr0qyOZIcBD2ThZ14gLcGWCjAL6l2BDp3HniVsmkdQPXjLp
SCVnPSUl79n7KS0vf8dutB3Vc8cSC4oHGlwX1hFq6G3ME/bW/JW7wxYxBbCrkaPZpsq3+is0509J
871ujMyfXlp9itauvyhT3klywlQEZ57UXTQX3xinzEmZjwQacMSFv/xWqRhJUmFtZCi5UQtAlzUK
FNaKn03ISLgMv1BkcGvDzl2HSNC6ff1uKtsHwTae4mp18Drj5ZQbXEGmdEnDIN6U1qySwSi9oDgX
RRhtKBGkKlTWGY/ra5aa7zZ10aMsx1ZJLdqQmpBAFSr9prunkQ0MYBPgdyUF9/kqEfWD6FJCHNAy
rWYY1WIkBJBhKcUlfVbCxCHqlV8vX9JowXJL6r4gNdN0Lzx30EsATr4CwDWWdm2ZxDCLnVQUWbkR
HFrOkFkj+5MFOtIoK0QllHPMFE6xRZetbfBzrFWQuEXvD2ac1M+2wssfRNsy1zb/CbZQ/6EPWK1N
5GuunVORu4moxYn8lSoxAVj7MVTGKJ6Qj7uPbCrvIyRXgX5hq14vgaBsFYVwjEp+a0YAO/5I7kCz
uyqzbqTpPhQ0plkIElKFce0Z+Q7+J0yVtYjJcKECplzTSuTF7lQ1fvO2hCe3OWuonRKt5pT6Fg0W
XY/WJuHK9YzYOjtC1H+/DDYd+fKAlWL2xYp8/hKZAYQJyslz++qGK1PlbXr/ERxF10l1g+DguRsE
JYNYnhMudvNlc/whIq7WozH8mMScccuP7d1ENL3FxUzqJrF0l2HqGy9dLzpE8PWl4s/E7vQ73KFw
4Qd4S5JFhe3nOnvu+Fxczrj7Qu2PfcqdaMRQvDbn5vw5W6yqdlhzHj72pitsQgJwLud5HpK4aQDG
LO5ZADnnt0HmKbqEKb0gu/mkugzHZzvZroTc97VqtblG20/5u7Ue8J3N4LmIl71wQ1pNGmNgkYfk
gXN21VeQfvG+foGmTL1s7EMFE7BjrWCcq/S28xNs0/AqoIq9npF8v06dlhkelRc9Jn94sdT9er7M
f285YfUorJyWNP0wpc8W658e5M+iJ53YaS7KP55hBjVzt69zemF8LOU6MY/mf3sVSLx1+oCKE6xZ
95w5sZ3hVVz8OeoFpNFVovYf4O+WABTIQopGT3tHNVDyTTRxBPyeiqi9MZvKoVsMOJXUTg76eOST
1JFFBs5p0+Rgge9TzBR3GyFEtDBmlOdVeuBsEs9Xgp0Cn2XpfIWOCbPu6xmNbn2eRNZxmrElfoXO
f7Du4EqdqKrqtPGs071CUPvyGTmkfIhox3o45vsqx7xp2wbIZMn3CTTDNn/do6rVtt/V2TA+feQX
5pwinaLswV0UiH9KH2HfZN5d+zscYU4vZFmSNLURP38rQtKqB94+Ul2QaT+kyNc9pFLkGgJIRuzF
oVZIBQ1tvQc8I/OyM+9Do9S+HPWE+q3Cj9yZnb63/VoVjE0M1lzM3TiWVq2oOlsDt06jVPH5OPPM
fEbb5+HjxMYGf53v24xm74NeexwCzd+nJEMKyABVfaqVqYJMI4k6ZAN/kQbTSwwtJeb33k8HvQBQ
Y2zswWZHDI6cIXqjF4FD5n8X5vssG2yYZdsNIyjRYLt3sjSoF9ftoALSp3iMQWvAey2HrKNicv4t
/2pfeBSbQhsCldptF7yKRCsmvQTOcnFtb1SJPCzhu1kgSBetntAZfZX0ywkMsCXn7Ew3mEH6bxSj
T2YoPJKenhgsdKMxdQVdyDuJSb4WcYUI+DlG7btxxHr/LsaZX7FWBVWCI7kqUEONdDFd+shjENvc
zDZCzCiVxD/sb+EsoYgxv7n0DVA6ZwZeU0OQf124ZeS6mt8A4YuK9WhUC07iXb3cE3Kw9X4RtFhK
VPQQvntZyx42uf1lFy2qlB1p+LSoUxdfBIOhrMFhmoG5WnJgY1gDp8GmOsp05FO3OPaCSEDmQe5g
TTu02vVHy3SY19HZR4BvyPMw5QAWvkU7LCd+BpjCO3N7j6FuheXDFa6LbmeauLVmut0J4RJxR0Mi
yhsfNVFzI7jqdY3HlrsQwZ7bei0wntpkSe09ggV/UYDnfaelvc3ncdxYLMT4EwbjlzVlek0J42fI
Dj4Av6+eafZs/PLRzKmRQmD9GAgyHPcHHkGapqaV8S+5JUDG5Z9LU+vjy4YgsJ4yLIGWCelv53Oi
UzF0gbBxY+LNGGXcZ4nF4vHFacD3Jf6Lf3gmnuZiBQQZ3DnuvMN5sECzRtx3k3CMReKmi3T54hW+
k7K9cI8rOkuePUCXTJDi/TRjqClOKuYW2o9HH4iDqsskShKOnvUHfo4tuzK+//T43Js/6YEIumjs
+9lUzm+4uCGK/po41MisvY1ozMz4+KJCHCu1h0qPKB96DaVQ17NBqxRlCLQ6HpX4yxzkgMIMuqjw
dBFJdpt8T73DXhMCy64zGiQUKobI+r+ggZuGmYLkniAZiUHYKMHasVDDc4I5s6EvtkTVdGN1Ra+o
bXg7+rtXvGEZmdtVhC3PhgJclyUQHpoqAeFZQPNz2REC6fhLDLUZUGG/n7SZpK0b+yMWDyhPXlPc
mT2agMAUFSK5b/gJI6Ipc4fgCwzSAh5Z9mrGrKheAfGFYU9DlyC8J8f+6tSIxWUNOyhbphiew7h9
4/tRfstuVmaiMrfivvr+pnt8WjqRzYrXT9XHV/3FCrecvNQqYBrJw6kWD6meHyS59UZ6j4LP7Twf
NwOd14hhkyCWxF2ivj+3x5DPexxsyoadb2LXYzZMkUB0FdDRPnua21anXaxANSfsShYgt/BsZ0qc
kIHp6fY6KMzmlDJUB967RcWYPVOWT6VkVDWGOGxivtXweBI/U4yDRZpu1g2caTYj2LzkbI2/xIPN
T/Xe2Y6p/ePJGvVoOIjIhn8L2e0pu7ASHI2LllAeHJxw+MVOO8guezJbMdp8bQn3SSwFssu0zW0o
T96dJfDhxkhfsDN94yrAwyj9zL7Fym22U7uuvj7PBlERQi9UvJdJqkh3/6uUSZcWtYLmXOgKmoI5
vhjvCZwWN2eaZfUCyFlz7lOU+rQMrCFH4qGn2jXhrGBUgxeVYGs+WNqk0pslkuimQoMhbTpxRE4h
jttQKnvJZ1O56FysrudzNSuQrqYhG0FWw/D7cDrVg2jF6m1hZy8ONGFeiqznxHHo5ISh46GZV2Fd
5yC4v+dK97iGe32W6+VIazoKp0eT858Mq34vnNzIRouJ5AHWp+YK7OJpuTO76r4+fgQSFg920qSC
7tx24st2Mw3YN/zBl16UO4EjKJQVJd2i/HJGrQwBxQVM7OUTemKsEGQN+tw4NGFiEiccY3ZOo+z6
CPpFwkD3VwKsjP96aPTlTRidlywhhKRA8pM+6YtKMECs/8MQ6pDrZCL/W5n3kSP+WYmaLDW1dCtd
1ZpTfZERDoXRsCwazvClRxPHVka+6eydWw+H7qy2Ko6ei6DwUL9w8cKHJxEfzcAUbSQUWGf5BfPL
RWwJV0ONHQJCGlChZm45m2sbrOQIHbbdAjC32J7o6v5X41DV+7sC/0YiH7aMVGIIxFixtss402T2
jn+CvetwDj/KncYeVH11NJMrRpwp3cRVzCXSEi1/UvyaJkn2xWIq8r6+U+FWR/hnI8Z6biMRD5j5
Z2Ik44hzz+fldT32lvesQ0Zf3ONYDOeS7paqcIofT3UCq1VK5aPSkiS2sxLRW8jiDiFtZSa01uKI
Jtiv7yrp0Oo+qRXFl1fKRYimP1ntVZ2Xp6ZUlWMHE5UAZ2VNhBFylk7c1utWXE2BqL88i2UUdW/G
iDzFT0rbAyKltvL3pcvKbE69Ga3w3/UwSWdcPPz86vaT8OMAr99PmblACnhcgOXbFZeH2TJUkoPB
2fMu1PYqS6M0PfMDeY3iAanzAKh4PGGUwCXDvI7B7G/Q2CKgCjNWa6VKFxY9jcLbhtU2/C168OVX
Tk1tUwdBA89RWhRIgCe7gQHJlBYE3IQhD/jUPVlGF40L+Or5MhDqS2vL5XiKAUnF/BrgL8w1U9xv
ORF9QNtuw+GhDUAeztECjIbSel2O4fg/C8Qwc23aCoJIVCFgURR6t+RJpeyEEQ6edaiuUPi5dOIF
WgR+73gznD4nR7ZnNsODmPUJIlchvZL99HkAkxJkvVXbYtb2NFmGEEz1poygpWKQ/SjgsINJxUKB
GHe5vidAVpr14d+0Q1RdstrWXMUgoey52fP1L/6Y56QAkoKCmJehPd8u2eILOWogVzWx4Ww/aKcs
YkUWGqQh2fQ8M7MtR+Bhi4+dMV/3ZXjqBZVOvBHHkoylWQdz8BCrbXZxR4cM1MFpwrZ/ZxxOGN8q
40nbdwVKd9PosadybUrFXDUz3jRY9Fqv4S91wr9PoTT12f2AtewEN4/XwC91VreG2y5U7OjvzLjc
LcqVgP+bO3Z6hqaP+RTqKogajYYW7nUpTPRQDn0RBAkaB1aNuPgKWYAx9PkXeHhpAICZdqKN5aBZ
lOFY8H3lS+v5Y+JUVxt8yZIqK9RHu0ABNdbXGWhkOb39TlC94uBAaB6AFCLypnoM7hnc+7UT0mdo
oERI0XvYDwyVT9zeIyyke0wYFfXzlarqGsVqSm4vUqigEOOQixseLTV6tBpS82dkqLMyiIc1EgQd
3RsJv/ar2LtrqkdHVEEJqcETqfSrfq3QvTcRH3aIlGUlkJHyMZLtHUm4iWs9RaOyD7+i2w3bj2L/
Ko/JBTONNS9TJLj9qhvMAb3LvyZg7DrGygtiG0s7JnFf7bMM7SATx2nZxFt/0N43vEiCgqcYDO1v
HoLGfCFXa29BTjJpZ611Oh7A3kA3+egGepTH3gEhAxu64kAX740QY9I6YUiYMkKiibSnxyXRGHCM
6XVdfmVlO8+cb2UU1P5DK4QQAh7075M6pP2cYNRbyucaC/FNjWmb4CW/VO9jX9r3Mi6Zm7wMobaG
4HP3qjjQSLXr/wLhL9+dRMYc0NqxJ6X4d7fi0rZ3tUKLKL+brX/KiTHjM3tffit8EH9/4TJgNoBq
UM21S7JZA5NXcOdF1W2bEmBeXXDRoeXXKfkRVwi/VFIQh/iaq2pzMqsoCml1JQzdeM6HaKOemyA8
DaFXVvtMKsi7tAQfXTXUUKuvNUxqaQNSZZPJOVKZjY6LhtiA3e9U8euHZJ/BXnK+7+6XJY3INpzc
vuTxaWjOSN3l3myxwYaEGF88pNlpdRGLZ7zZSnyD6ltqeF8QL1TUr0JGB1nWB8KICzZLZtLrpY5l
a/ipNPKHqWgsSkQ7DRmXfcHFf0B+tJSkm7/8w26WuAGifSq2qA/KxPKwMJe/KSflb0LKU1lOFzry
PSiS0irK151pViugKqYlQbgMaK2pPGiQcGi8fdTEi65Vf8t0tUa2esKGSEHgw+agtzKBNFU2N9vF
RAkptRnKnUr0q+oP/IOG31e4PK343t4jXD6LRk2pQEP3iwvm4dTbByHIs/Cctlb14IQgLpEKNwWg
sL22vSGZZLBbqqjJwjv4UJfnCLlwd/HZVsV/5PsJTQOYwPhI08vfRu+cqJXTGV7ZQuEdDYVTW/mT
JM9Ou53cLqL+Cut0gqj+CgbAcnjdGRaRpst2yW9VHRU7v19HS39SHcK/JA6pPQG/qP83oU2jFxYp
yil6WRPy0hL/LpoCST8rs39NnVrCAQZkN2iYT27sjEPpgfh/DMFeOctBZXRGxw8Tq9MUimNo/WRt
0ye5yyqOncwPFnTon5f5q/CNup6ctuSebSkfHA4B2z6FO4t/+ZqlwMo9GSsFFMhgKlE/piOUCeSk
Op1nWjtyL+O1Ao+IhDJKUGuJrs5b29uXUenEp2ke+H2d2/kxNCM8hCL9X/VQagIQrForUlO01MyA
vuTtCFyKH/lgdn3DiLbIWvKuO61MFUiE5tZhON0V2UpkQojhPjjX2o4/pCJR2X+vhWig4GMh0J0a
qa/U5hCAlEevsvjm/AZm02xmT2p6QP6sAxmuWhSNaf5LGe8ZV1c088sWRmIyD1OANRYx8WGyurC8
cTN1yzGXc7/3rsgqMVa5d9UnvPM46AHYSCoSLiLGiwjL3pY/wsWNxahxp4Ck0UR5mHwBiqHFsp+A
wpMsi4/dylUKTpD2hI97P9yWYnEad4jJ+zXOlPHR3MmYq/rLZBwzHzD4tLRFaVpS7OaAKHZRi+Pl
5P5OQv1wHCYVb5Xhc5KHslTMl0kBp44zXq+0ok1ZhHJKhbQhVqCnmixtR55DHBbNVHT9URXDwlRX
ksjvMJUEF6kpG5cDNDTOgUtvqwIOOvSiIs99LzHyk+Q50SYSKhBGzyNfK/DJToHeJvzqPF9x0cu9
85zTlTMI5YTsGoC+V949PUl7oQqOEdiYBiyrUPIlGLnS4VXYNNUK/o+1GXPiGlWHjeKVWNWHfHFN
L4F5hJYQT6G1goVCM39itlfABGjl3gkatto1rI64vzP8vYyUhwpIvGVKh6qTx/Wo5GmEGw4yzWiL
MSXcm18u317CDz+kml7/3FFnqteA6cDRZjewWfnj3wwbmBd0v/3I/94oqxIMbs57Rj8vA4D6gaax
FbL1qQRvdfx41k5Wxlw0UqLxrLJN9C2lMHcgmG5wBQf0ElCvpJaEU0yyRPWCawD2GqEEU+csjccT
KWGK9kquUFtV+XNgzZdQ81Wkiz4z3AYU3jxBMmjMtSPJLzAJBcQPwqWPpRrH4CLbA2Tn2OVU4Z+W
Trnz9ZGllbghWxEdrCdwRExOLVKHhqwpQyPvi69IJNMhQHdu4FmFQXZotMCCb4XyimANA2M+SZjY
zJ0Ly+rqMF0U2q0gu6ZLWGJOFD5RZWCMyU7wFpwOmj2SvwmJYTKhaFiH9QGslcpdaxJRnAchad7M
jNgN3VG+KrRLw+TUtG6b+UT4WWL3Ho5f87BcSRHNcQBBtz1xKlBqnXFJcevbsY9pKUWz5kfqKvPn
X+Ad9ir9yRt/17+iZh2P/p6VYjOF9tj8pFf+UA5I54L6bKTN3I7ddgspMdlCtrCJMKeAfChYQ46d
Y+iPJ4jLksfBWDd/mufS2WhWDsFEbUN7PI9YL6EDlTvKnLJyPFyYSFU0Mi6bPxJObvF1EEOFcg9Q
fig+FcfKv06Se0kD1ZPzCLoYS5krtw6CCVdtI2si1ueKJi4nrlhpOPN2oFXFlR7nm0Q2iWOY+t/u
4QB2C1vw4i1k1P5cdQQEKzBOE/jw9BAJatP/sVdxOulJXv2enO3pBh/76fU2PAsWY07QjyIEIndC
7lNkwe5tBhWp4m9A5VLac4T24jYsK2AcSHebM3NPgGLHjScqkjfbyyhr3Xqz9KqAfLAdViNretW3
qBt7etjrublMw7OsI4ZIxLUySH8eLU/8L6DTE7UiJF+bGnLklQeTujlE0FG0dDbf9ZVlrQZ9Izl7
pvAHbBk3a7DwO911ERSpMqh8ILAUIsrg2Z4zxd7kDFPG5aSR5PqmaybcUQycmi4WqYOF4f3kojEt
GiTZAjfDKB6VWZqQs1Qh7ptST3wZqy7Du9eLDwfL7r+73ZXId0//mxliApXLhwUHcMcES/KxxSw2
u/wS8Nvp7zidgAZPQXFGc7Tlw7luw+xWtpiAsBDy5/6MS1V6nsNM4L7kjB6L5XsnSObWqMJfXPG1
WcD562wiCnpSoxrEJcIgJ3OgdPQURbycvAroZOpEk0HhIoBa9zrKjlyzrEttWiu7/7367ss8Gi9u
VMVzrqv1b7YmjL4xK8hsGIU/tT0t1fQ1iGLO+EtD1jTGhSV9pkIp6jm3vj8dj/HLVISfxxCW8SV9
QElG2IWOsthPM1Pqf1uJtff69BRD4ftYix+ppchraT/k6SsGQ/XleuuCYCWSD9obR+vGmA35kfFg
KyE79KprfOvzvQjo4PCxFtrrVyo/V66VGnsYJwlhL8RBfuqd97LRuWItCummRjgkqrC8xx8Zp8+2
beHYaAkmOYsM75iTJNacsmHLDL07pl+p5q6+ViS1rjJWfn1TL5G7MDfT+oym6RG8I3pfk0i52Irz
ZnuscMxzaxnDxc2FCTZGRYp3sB7fdccWWkiVDAuEcXE7Ou8HGW99kUGz/qKw5iDWTyjXf8xl+tHU
cmKU4Q5vMQ/BA2k7A55UVoYgAYGoBmBxjsOhawM+Hkfh61H0qt0Eg4YWC8oSyW5SSZIIenRtAJjx
4Daj55zRIwJIu/4OF9SLAukxNFtxNg3t74HZ6+0ZcdNrni7SWfROdVK9Wrx+Yee2vHqwh1xWDjH5
t3iBngnKsfYUByMcuAYlJOaVJydaSL7reogsYcBoBzM0LKwRRDq0fwu63E+qu89Fk45FYhKOdrr8
T2ESFXFWGJptpUylRMgC+tOIsbUGHlsBr/q8qLsBRsGhTVLHULTzVaj8/GizIavWIjJ584HVevaC
HGmPq6UmRzXdUUGi/Qs2k7IgyKgGm9U8BFrrKBBBBpoFQ/030wkgkBjX7PN4sRtHbtan6S9FWDdx
1xhDqvi2oNQhCRssEeX3hz20B4G4ga/Yg/oHehSQf4Yqt68dsv/17BeEXymmVjLmW3J8oOncax/x
doceXgKw4UtGZ7649TrguvrgDlyvAa+5AKi8G0tYnC2a/NufzjKlHv8o78q3jDsNDp5CCt3a3wqM
yVRzVDgyT0bDuzpiiA1KlUd9VQlf6lm62LgjwX/bTahR9UQB0KYZp7VPBzL9TURAUKBFEmmzyPkH
7ocgstibLHiJEgZ/BXYsfpCY5R4ah1BmRrUIfx9i9AICgJyzQW22q9459wxLzPdsLIBRnr+l6GUj
R9U/Q1TaN4Nx+Dz1hS3SLu/Kbrz9L6RX8vnVbIXcbGTMU0dtL9edV35KQXUW3mEn+ZjslzxpMfHy
+GabsRcle6CQcHvxlo9RFGxc9SKfoJ5kATdwhVDiXJgoF0trOBRMHjjTjwj0g6p3SJnR2kNAr++D
6M9sTACmGqcxsxFXwO8YQ3QN5o73KpBUU2N2UR3a5K23UBpAAYEolT/LlxRVsdQWWYcon0+Tvb/m
XCb9L7fTeuaCZxOoGLUjgyUc0AKWSlyRM8eqsRnGhS05fFFEDKnni55sUTfj2e+tOxQ6tjLI/k73
U7cwQr3bos4MSEayG2KSylRyLDkX3uFILyQ6ONn+rBgQlqULQ7zJnLq3Vl76bAWKokS7+cNNmzjs
DLeIZvLfEw3f9kqhEr+Onpht8NwxBkWEJwgBfPiSsf6kroU60CY8QlP2wqGYVik3oCaqTmpMrEYs
o5GWeTGDCMvCwR+AhX6u50LupyWWyGQb7ooFqCkXp7/+7Et55mUPEnDcQi1f8+TOFc0ryPo+gE+e
Hk1wLABACfEh/HiDV/Vo8MRgyBJwHvo7pPznf+sKul2Rh0lNni1/NjRh7ovMbJ8hGPhQRh8KG+eL
bAGLjdSYp254kqVG+YfqOfcZddo47mi5CiZRXaxL+K96aG8RnmI46bXDLA0adSzAIRZumCfl4aIk
EyhuzxlvBwbUcY97W63iPxetxuEyIhOwVMxNzQ/waYf2H8fj/bM4qjBy5+jFepMYR6h4TVp4lODO
1XTndOG8T7yw5RvnQ6e06bHS1g9Mw8VqWVSEvz8/Uy8gCF6cPF3OGcR53u9l3v7JGouTY7kgwwn4
MleFsX2g34VYzAAVabQwfn55viA+IN6HiBaunK9vQfe4t82WcTEDuLGYfZ+7itasxDtDEFBUHVHi
Quzd8E2GkhWVt9U5iWNIRvzST6FfvIg41yCWZulVJeM8As1UOWMowE5DVDf67KvKo/wTgK/N815L
pscG6XLOQbwyhaz7A/v2PnMZ6Z3UVKWL/IKzrpP1SzEad0z3pxJVCc9x7rd+jI8unb53FiqNhhgX
e/kn/88P6aJT4JF0YSf4hYrWD0XbX+hrtoM2o4bquq7E/D8bIQ22kx870kOKyU6FHcFJWUg7U8n2
42KnNNA233bPZmAxj/a26q+NJOsFFxsCjn8x9fr2KeORWV5vw/wAQo8gSh5ChRWZSsBYL6sy3SzF
Cy44BSq5rwKAEPBh/LM8F4lk12y2Vb/f4GC0JZoGoSjIR91LiSfxWCwEvH/S0qjDv3b5DhNnAEf0
n/dpXYQC/e4PX/WydrPxMNsz7stwT1JlKw9oeU4TrzeN/FnwG/todGkXmMIS6eFwVxhz8BlOFvf9
tiwg6L38VLBt34AXIGNPy0drBuPTgdCgi6iCN8hCR3hwT5lSN9mL0VbewQa/WD3qMfmOfPVTNqiP
VQZcebpqbPdj1BYX7lqS6rU0YmZ30/pBxMb6cl8XQWnirLdkvAtEX6vPNQ/UPv/9LaTEl9Aaz8jO
B+CzoMUEIhLbwBpn7DzhzFP7otsxFHf848pmNgV3Io6d+KHxQUYjxsmOUxKkjyXfs762pksJIjUx
ma6g/T8NCfm+avDbK0VjLxSbKcr8GNlmgaDt3cJPbSreKC7MVTt6BUFu1uweG8VB10v/jIvtM7+7
ItDM8QBuFfZGze4THo4yVTzyA22YwQ40hzUtONpUtFhSbsfTaUjn+eSjlnjRfA2AEkvn8Anri26p
q6xaS2osOQSChz8Qm+USeo8LWuGhnloLay2FnHxwUF95bs0v/XXVnHcfMIvCgQhN4QO1EzMDZ2EN
hO9B37F+LVK42OZOLOnjL4wDh8/z0pc52n+dH1pgBEjCkanCTdxBlQnhRcFoyYKxTzBqJ3KQxxOJ
0eEOB6JDhaHehsZNeZnV1s+/lWpo66KzjQKEwwnEV9dleU6YFvGlsSY+zr8JbGC4aLiGyUVvigUA
sppttWEK5tmsk8oLu8T/2iHMSxvvjllg9f7DYRNJRAjUhFuGWQG3EfCxzIO7BjiUgi1DewJ1GwFz
AQX3+BhwocJrdYHH350f9lYQ3aHVYVY+rmwmLFvFkeFU4KT+gMo3ndaDlONl6pRIevt/uR7/GaUo
56YM/TPkF9n31iHcXdY135te4Pb+o4nqQ6bkmWzDQELE8lymWkJzg1ERVo4AsDAekMJf3efITv1R
aDP02cE5QcJs4f/gU41Dc5CfbQA+1Jh19TzTZnxmjSxNE+kOJSG+swxiB3g6d1E8n9VysB7/s/Xf
27TVwvlwY45veZ1lJm81PY8BylNzMhQWFCVnPRhYz+fuaZL/UPwXyHIY+dhzV9js0mAmJoNuYM6W
IhK/jiyH/pz4jURDliTd89gGL2wgHNpYKR8xxFGKowP7Ued3cSkunsNbFM5SV5MmBMChPfVBmfm+
sxtha3zbhs0X4iWzEEDy6hGKJmhkjvzxwyNO/Vx443P3cC8C1jHcnCB5tiqyfFJjUevL4dvMlcpO
5e0EQ9lOH2BpwCi/E6wbuojQUGqmB+UFBLYc4hrcROPSN5rbwSjIx/IUse6o2jg1sZEmXm7DFBm2
ZcbMXBR2sRsnEz2tpEQwF0ChrMA/JninXSWZPhTF7D+o4ysaK4Sy6AHmt4FJKQcAXdWZkrMVY3Ho
h82Oz0/Ao+KMH2vut/4MbS9l3Sk7Kcjt1g+aa9yX0tPy2kQjARpP70rM8PzK0QE2lNAvF7Ob7wHV
fshTxKJESVwe4seA5EqpoG8VAzK/xvRhPrEwtkZhmQlxxdsNaCL3NHViRUFykTtWeItXw2gpty0q
i5A+vpecHgOicSc84Zy0PV001ofaFjlg1TVc6RF59dT50r0+ANvDQ32M3M7KM+Wp0g3peGEW7hZR
l3Ik963Ece0S9Dmu3vdpabNTUFFVlKkuoLp2aIy6tGm2VyPE06Dd503gjHXRbQneqR/ikq3MTh/J
bm5knGOlYJ93IUTh6amYJAw1GEbhE9RxdIzNrQQQcQHD9lDBmhRv7FJqkBGka7jgT4JAQ0soMIKQ
5Ngpvdd+TribwzwahgrF7OtLpSwmbiitl2MlQC7KUE8XHIaKJwtomHLqLKEcXGnVoCIUF2jD0IHf
1Zz08vh/y2rz9UMt9I03AvHbN+dx9Uno4K5CtHCrpdi1cQkxCelwknDNnwTjdph0S7gKycq0rU11
eQdS26H6H3GGoeYxJeQtpANM5zaazNjJrxJoDdU2Qy6c0lJYBhtdrtuTQJ7RGLohHf2yix9gTp+r
S7yHYtbj4Co+g5gn2Zit/qhqv7y2ZzgIvD7lgPzD6iHy2L4zdqHfStUQ8AxIl3NPS/r7UaLwB78z
2kgew64TvtLJ7/7BGfRYpA8SxNrXAxsPDbGIvEg0TedEuelTnxa6rs+kk543AZnqTt5x++A/qhwC
E+6fYc81eG9TeZJBsIvmKEwIFTYEU+UIg6CP7b8bINvywmyKTNiOO65ep283Pxe6dE1ZhOrdpd4G
gDctiWf/cTZx/UOtisMNGjh5uYb8AEI5Eb5606UuN/2CMyGwXuBQJ6CFBxi+8VJSRwsTaGHzRrRB
5YQPYEBFP2NTKzVAXowJoU/fqS6o+RiqhIzpsGoWOp2aBGAwGG96MzYVIGgMOIu+/gfrxJKOIFJA
jbkQWwJ9yZpqBe7vKDr59ZgHPq7Q3lUYeJEAQfLdQV7NXYQIDDSrK9Kn/0kSqKVxWGDN8KM6ymAx
vXKoaBrLXkSicbRkk0yXjSn1NZ0TcD8ac26pJVWqwNkUpssMp7rutIJ/4m5ke+LIcGpykbM9rhhS
QaZZyGAn0DiFHVfTrnXpQFFHe0scH682m3pr2u3fNi2f9AZcdevA6TlyXWKAk4b0q+ZqW2ZW+XkW
Z9fHPq5cnjQnfZlwUUGL3GJmMy8nhDN/xTUr4NlTvi5WZIy1nCJP4u/pJ1FgqU2Cd7UYhpCtX4m8
PvR82sTYcpf+ZOKPgGD3RdjHUvmAC3P+i+NJ61Wp5scA/xW1II5H3V1SrLv5gWrN3CZA7oNfiThM
Y3q2dO2SW7riguycAon5+CA0sSqIg+KUjUfVJY8QcvdQJriesUuMX9jSfy1WZOogzGuQmx/yVVo5
lrBUxDsWg3F3ZhxrABm1uaG4zNNagPv4/6+SbW0c/8lV0Jvy3qV+EMOWeGWl5ZB8cZh/9bGn2qDv
f+/yzRA/K47bFdmZi4YM8FLX6tFuWIlJWYFjDJnwl9XGbxa7Q23QpL4+U6P5nzIfWsx7W1rI6dPK
T9CXZ8b8S122vai9a3Qjn7QdAOKp6iRTBJflqUmv8gDTzGCZNkrTBYmcddgSlGuNMmvV0fyVjHx4
l3r8SjsXsuC6oFrRYhMwmq0ZZ8yRv6GMEme0EBFLodhMI05+oAu/5h+QtQzIShesQpWJOT7cHRC9
/WeH7y7FeI5KEyERUsliZUHbOn9I3q0hOgYCo2DATRK+MddTLMJrZrn7/ChtGk+zCLSEOwbpFUXx
A+HR9QcWJiLoRd4dQjvO8NRnYKr8EErQ8HzCR9uxEk6enicUpfQ6s5yfEqWNOHbWo28gOO690ocT
CNOfsBMEEC45M+pMYhjLw9P72zY1y2Xh8DFOICa6tchubMebzoQhQGulnxkrTsQqSvcreRUwQuFQ
DMNVtGXywkRSjb1GFxHTozwmj7f3yXsRkmd9TbN+dTT0GhxNtCKefLE8jLorwhTP+qJIRZhrCDYh
v0ShpOEcxMBIPDh0yfzNtcW0RoaD1t32Wa+BYa2iUUNdPo/jhCg7tZkoZX5XGOio8wkMD7B+tsHi
BR6kBvzlNjiidPjmc76+ews9jpery2m++LSSWlRduH9U/fP44ZPoKcABOPl3W0Kj2ygdn7ZNOEp0
dAU4++Mc5emBA2UzyHYhHFgZFTeVB9gRbOsEwG3gilnm0v87tlEXpwt0EYU7wDFpb8zDEwNRhnlq
6ZQrrt7+fplFRx7J0DXnm9uU4h03t8ZqgePKnV/HuQGbxtgPLaRdzniYY/BKC4Oul/+coK1bp9wJ
8ayY9DsK06zOARm3YOdZiuJ+tsc0CCq/KxGFUc8/p0p9mo8NYNNSEpkUqWHmNp/hexYODPE1bvyA
f6nH7gKULRaS+8RhwKUMNe0S3VqyFiP+TPzkXldKqExul2zZxaPu/F4nuQHdIPPwIeww5WTLmDwg
i4t7fcHwmttxsrCq9bp6rbS1aijLAyKyxARh3oncHPu0nT0MTetE8A7xA0VqPFe1zbtoIeK+Drew
SkBc+VcbM7/4BD+wiUNMfOlNynSL+M/gXtfPm1IqiGVUJ+L3N09/uKuGsdWIGkUcMsuRjc1KbOD4
/EyT9vEypWYsX/ozBtSeAvgi1SVrLJb6/ya997aI6exq0ebkNwRrMrfhpy0yBc4iAjVcuq1/4cSl
5L3hs5+JuaWtfzMsrG8UD/Uy2hShnO0xq/L7zThak1MLKlGvVQKDmZ+h4Wb5ZA4iGRZM4SlHuSVa
WMNDsPnsNlXFrClhxuwPTXH6aJOXrvcXQUZnxDa+Nc/UVZ5HsxYY+tIITfWw/cT2vuLWwrXtTqXQ
t1T9A5jTg3rDdzZ57pwGK1C9sWn1B24hh6nGCokdleso4Q0r6zk+uW8aV6lJXB0eN2FTo36Lxfzy
Vp0pYR05XIaHTIPpG4XtbrzKyVNgbQwHZiSZhLZDwEYZAyy331XWktQk0BCXr6ISa+Jhr37A8ea2
yBdVbUiSHrmOlSqB0LkuqJK26hMYhOdW1fbawJzyOMZlxiM6u+A7bsKKlKG3ai6En+X87qpJQcB7
9tgfXS8YEeIS0dru+TEyGvtT2ZICyEStzoyX84T7qWlmwktBDzL62Y+pFePydzhnJMPHZL4zUdt+
FzUTz7PW++gFBkT3ZdJl4Ab2QNyIDiKg7tz75WVjLK8HlD+sL12uwXRrvnYYoBrB3ZjCBzBSCRQA
qTvD5GQWDxh5IeDzFLZETYCH6lvF1ErIxVCN4YXxtgtUKyK963JnzsIEzeo2yTp38w8KvAjsLeaC
ebB9TwushTKzeHv3Swppz6GEkKniOQonijRCoqLhBz9lo5RTCtATsIJSVuackiZIK51A1ENeFyMS
Ow35alEbbLN+aAQya8/OSmDhBbWXLz2NCHIik+MLdRXmgMjlbFDpAs+7RUQ+U1B3o8CdsYl3lIrs
7+NOzr8OSDNf7h/LYoiTLh532QsnSzXV5vIyKP3PA+odClVVgbLfVht/XLsuAoIyqCVWv5v8Q1SC
YzFVkWcOdiKH7eTStf5K0F6tC4wZALv0YLz4xxDbkHPv6zcS/3IB7t5dTuifq9I3NqfQej+YIQSa
r/R4XC86/Jxtss7pTL5QXoW5QVa0LgbQfPjYdobz2TffqKNCiIJxjU/7IKe+/2n+phDsZdkXlsmp
T86K5hGjfkaLcCzwK1dwWhPxal8sAV94v1wc1nGgFE52h+e79gz+ZWgMqd22oTrXt6TcX9U0dgRg
yBanb3mKqapReNEUd73dgjCd3Hl3+avbPhwapnV0eQK0jdo8arkyvweq6KqT/qAivawFnmCbNsAM
s04n6+9wqQT+Yr4KBEnu3tAPI5dkyWQu8kjwerfbcacDn3OuomKaSuCNCzlPQ+rWfxfRiZ8Blxj6
z7YTP8IkdN/WW/CrFW9/yo9tY7X3ABdpua+yHriCx2jpTxhGdVemgV9XOM8XckGDEeDg1z1OV0sy
qGCCHMZdX8mWRcvFL7gcg7jkTNsyHiOOfBj1ClPJi4dvh23ta+KpoOsPBNQ4B4eWKBPfSPr/0iBZ
YI3IpSlBrBJSyI4ptXRou0g1YsdJvEaG4gsi2aMyyKIGcQ8FgEe+6fRZf3Pbtmh2LOIV3hL2WblO
taoOKUtrfcr0Cb2RytKzsoXnZ4oZMJRxLYn3HarGgT48UF9DD6XHKuNc2AjG7Z92n8MCzBlgzItw
U4r2210ugyVNUr/y3oD3hlSYAHHGbYXClOeD+WEFtchkp9/GxSgBOzh2UvKyRzLhbAu62eCfjm4V
3sKeSnDkxK9Pd/JDJ9i4DR6CCtLvSiY3BVMR5zg9sM/7arwJFhututtqbblz/F1Ndg/lVRi75bHC
Ur78SqRSwu0qq9+menflbcV8gsLwc8ZsF1ozGlUVXlVFpolpn7rxNUMXP3X4JTTR6IUD0TWaTUbn
IQ5iCFJTAyQv24tG0zj6yc4fbuIJ8RP0Cqzp+chUFJ0EJKus04RS4o4eGhrLxfKEW/7eyH2G6FkB
3ueyRq/OmSqOLLD8sA3G0IMu/ZthEDYQDwh652d3NH2yN+TyTOYgbEVk3TpuxXrGiHOjYbLcC0k3
5Ig63IT/WjL0cbvX/IniWEF9qdZ+TinSAYO6dHs8VydRpXFGabdu7MQX5NzEQ6LE447NfPvhvQ8Q
2dfVQKhvej6GqNqR08olpgXWtzw4JMBN4dumocUay1fRBQW8hFq8RHTcFhR+r09LWGYNazFCUGNu
wLdrzBFMcKYB3duUwYeTPrQSEWfsKRgsxSg46JVYYfur4hFgoFYLVW1jlwxQBRL+X774dQqLBkC9
lV+I5mfTekhh3BSH5UhOuPs3QB7vV3hduM4zv/5VxP2FptG5hqkFVc/yNNI5quLj4qoR00FUhVyx
p3EV2PlC4agpkXeZNSKLa2YbAsRoB4AuIo2PhwYrPHwPrdeqDEPVPZ8W7vjrFjC9vT2sKwVAbiN2
I6gswc+LLybnmiuDkNS6kSYunLAVfbQCRUvPIxEFCS0oymnchK2iguo+0h4HoJLV0G1LE0EKGZWd
XwSWGTUUByXlg+VQiYsAw2BNMQvIU6IyxF+DzWBlliZ32Q6NBLRftE3svbJO4e6yMAeW7z2MkY4/
YmioDmlh8fOaufah4Z9QCS9ty+2RQ7vONtXGoXjGsJD6sjFCI3CYADwBHLp2z7GAOOjUS/rnprAi
GeXEQfNDe3qW1xRgLNU6UmGnB+yX2UhVItNg3zl3R4EjPbHriJWEzqk2Y5+TzfhyqEu9yaA1+ySM
5hthHZ+zSA0OTbO8qD5ocuXXIA0UmhI131mJck+3ietAeu3EejIPPeIPD4HVpZZeVvauQAwmx52j
CpeIz1PZ1PbVcGF2CrOncnQMK/tzfLtp80YFUIUzQERZK59r48Tu1ZQqdZAf82Q0Ple9KaiaoJ9t
1ChTg9fsv5gtpYvmwxHY7XaAbTkwWkzXm1S+4g4qo2eVskYhGHGSxziuVzWiALgQ1FO9mCZ0ccin
Yvjt3BE1aWg5YUV/yTqK5qrjkqbDIeeGFdDQg7jvKdZXIbTqv0L0mDe9Lgi836WwM7uqZsvtzHTt
nPo3Tjp/wa3GQkhrOKwSjsjLgKSrEBJbGMdWyELbznMYO/eK5pbKFgGyl1yz63aEXoO3MO1msVbS
Rzl9x/a5qNscGtogQPVR6SZQEeyCToRDvWUAx2eQN31YHbPr2LNPV22xyMADXpg7mqUmSsjrMIUl
PEAJ0DcXR8OEjFalMxLf8ZB4f1uIm1j5VgktaxVdB4Q54JDZkSnNxS6SfLijB07Znzj+/K3hgtLu
LfLFXalCjPdhY1Zsjx5zUiywEPAD8uw3yXBYQCBxGd06SnK1aZsAiNobV+jQwCRZdM40ZP3b5nrt
HR8eP++R1MBIXXE+snUFV2lCPanUl7pDUA/M373d0hgyHkjp31HYP8g4PaloaUKLE3qizAl4XxZ+
n03BKkMWgJIgmqhZNwjBuz6aauXsa5BolanXVYbKeMhFaJQLmdI/yuxM3wt0an3NiBnpwpIsK1sx
BJmci/GB5QHhcTlmiByAkZhegFgHqa4VYwRtousjt+3dyGJH49QYNLfGw0cvY9qT0B+q6t0hb0ch
77IJvjHuqcxukq96yeukFiudNt0APN6CkvwKixBZrh1KK9N0iLAOUm4ApF6/2PqX97PQFkZ5+5Tl
3hq+USdP3uJ/e+nKjDNw/mbEnSV9y0YSOby/o2CC2KBBEc8YgaI1jNIhrG4f52UGDUGLm7MiNlbm
F/iCPQwD5kdKLdS6F6SJhyY8DJTPQV+hDyl4JXy/Vl9tQ2Oqnp0p+kfPE1PlHudewUTPRc6E7aBu
ELE+dSTXpGbD/FXUxXtxwg3U2lThsp5LwGoSsrgOn8pl/AtKPh8yo2q24Ceb0Vk8yaFh41ZoUM2m
yuCOAU5JUayD08sANKNW13RQUwPfzYa1hYF9fips+xyax7rdUL0J/OPxPfqCpbJ88Pb7yHZEJrmU
qGd4++GUW0rAztWXl8UoLEIyRDVd8R+v9lfFJdt0k+hfAn2S7JXE3Xy7NuzC8gPQKJ7qLrxV2sGw
xn3zI7B0Dav1pxjdyVTFBKRC33W7Zqo+hF+N+hxaQHh2l9/v8dD9gjtWYHoX3nIDX3xQUpm2R1A3
WHwWpim+QdQGOuBkMGvRhhIkUxHU4ux0P2mfCjhxAeOBNOFioMIiN6nQtLxqkfPRl43f/3s6t1yT
FPP9391RWSmFlXLSAL5Upvma7pZPG6QJ/riQdNm+ghg9gRTzqv2A23qIwtpGK1uxf4UDyYqkIw7x
LSmlejuGvXu+vgudn7cblcLGdJsz31dSXMP0ufrUKj3twyXCZJJoGWwyHNKFzwcLMMdegJFCamtu
YKatqpfiiqX6cCRd2PM+lzyCcIn6NF585RoZPvz83bsHFAkRrYEl13sFe3w46GVEgWZWttbl4rMF
L84IPJttvDA9Ak0369+DAjBR1eOdCD7NlYOtqs5R4FgRZvRaaCc8NGIwqC+cqa5aDH7v8TZz9tv1
TcjUXDbYVVcK3F8cDtAKfsil4I6Pc92WJ2aSG1HnY/OycRYm2P1SsMIxRWi8JKTGuB3K5w7hqpcs
UO6Gwot36d11jZr8u01ZknpmPsLYKJj305trFfPdVOD2bjDu+EaFXT9GwDRBV9Tm4X3leLyjo8/I
tX8+0sSerqWiXfzyP5suN16h2WTb6Blmjh3w4WWXoSSHuL74HeY//HmQjYWYBk6AyHd8wq91/rnX
kn+V0gYglT5vKuiht5eTJuZx2kxL+UsQnPmRxJiF+N/CgKutxgQxfjZ1QJwojKzQ/3ifKjYaIMxd
/Hx81uYmAsn0oZGYNWgeI3XkcjzY0tD5+KGOIZIsqhLRJ4KwJwXBzQWXi+ko0+OXv1LWOH4k5y0G
39skhzBlfhKW3kGMuns8KpYJZmngbxgiskcwc8R+/QkGuAQ1uwlkteCqPi2TF0am4J1yjF+iWbMv
i/0gzooUCwqmkCZTneMjZPRKvlw3l6K0v3iLNPDyLzqw+sZaamNN+lO2DGROBa9MIR6Bp3xoa2Pu
1bJTPfA7nmFfrml2qF1x+7Ur0eyZU3KtatKcoFGa9VsnyXttRiKcSeE5m0l+iGxnKDfyMidVjPTC
Tv1EgEXwL09fp7Lf+aGlCbU/67zlosoHc8ET0h6ztFBLcUFOSflD7xTHO0lJYkI9la5NoasW8y8J
ZZvZMzsCrGblAE8n/3cdhtoCfjeOFJnXo2eSpmh92XujC2XRJ8KolZt8S2rA6szFpgmDUriA50vk
FldmF1Z7xPyAQkBK1m5lc0EYGm6I2cW+CdizTfA/UuQs8ZtifGd7QhMfFuO3mLOCK5xUHdm45R6+
kTk/TvIhtKfzeIZb+k762+YuzvxPpQ4y6oihjYsuLBZAWVMDt4OQxgYgp1fRgZ3pe1FLutZRdsat
JofCqHfWWbYHdboxemEnoPKj+fwnwWDsYRwdqJOwS5kouf0HiAQ07zqZudZMlADCpyuTGKuOLxsi
Qcc2X83ENADag1MZCMNs79IZqS1lOrMWW2JvWrUlUlTCoJvwPneFAC6HXbib70Jr21Fzgp1OXQCN
0iUCkZdyvsmDU0MK0Ynd6wSuJfqinNwlVir/6dXpan0HJKE0XF9CUv4CYfh2WCIgZ6nuTRX9qUOb
wmUj1lnGpkpp0qFuhQ47kv/+pK+Qe28/b6ZTfZaf4ZcNqC+AKojN4QIkgUh3DZdHJ8/7p2MYR479
jzXAXUO7RJYkx5sQ0+m8m8KPHfOxDFxSya0zDP9XeFpjH51CBGH9SiOQ9YFYnF8l24U+73nm3NhW
eDEWGId8ptvzBZz9onCYRQYe4XxaIzyjMF4nsMmLDZKIgN1jEnjtYGms8dd5KCK9nJax2whfzO4w
NoL0komvLdu2H6GEFNBOQD2GVMDRMII7vWzacP/tQ93AwNgh0HuTmUkUwP9WmPXlY/xPL5WHQhJO
EwIjAiAjkjkyVjRiDeUZ6tzcg1NNOCAt/LX0sm7kl4dCzPnFVvC75GZSbER0Lhi21hCdjTb92Z7e
1NFdSmQRMjtYagzAOffmxKUPI8ar5rI/H7gKGWb281TTFz1T02BTt33+DxSZBdZ2Dzfuxlp4CXfM
MTrb1z8IIDOneKNlbKC9Va4owPfc2e0ND7Xj8IF2QCGv4IeykMGFw3BTJ3v2xp/bqiHfGa8c+TRh
+Wklkkv+zXhctLnkYUTz/3x2IYsszHz+phxyrSy+QXKuZ2wrxhKiUKWuP46jUndf2vvTFimt0ltT
b53f67FHe/hBjpgBXjUBJYHCZf+Kdpe8LT/d7DyGmvtukxPad8ll1b6aKtZlAy8OIgP5xVD3DyI3
Yg8ejTpvoqqke/a6QkiKeKm3bFwDmCixHHhcdztDRlyDaa5QYF5Z9ZIw6dal/ugW1Tvk4yQIpugo
BcAQzp7KLLxgQtaA6KPTLV09NynHRuDhYHVIVsnQzpjR5JNmBXkc8pAOWLTqTMMfZIvyv5lWFUOX
bnW24Hj8PuTxqnq2UDm/Se6zVr1tFqtPigv9NmEng2I7i4vwujkNJzmF7NZf4sCWE/7xKBdar4rE
dZSzWLs/4MtE8e138eYKazSsubknl5+ECreYxdFF+3H0bFIU2ObWixLwIORxJoA1J4i3+Q0SZVH7
EuaZsPYBgt3BNJ2Mo2Wn8obTo4rml8YPlb/grWDrQqTo23MmrM1W+SllfrLTRywzXNhxXCipDe2A
LFzV+9N42Z6Trl7AF2gdFxSH8ar3R4bZFVU9ehJoot6+KIi5W5groLfE48oDUratTkmtZCNDPAV4
SbhBG3m2JoEY5efZJEi1UWnkw1sZYzselEAnXJTmuQ6+Quyjp+GbyGi6oMDoKfmvctqJJPhX7PxJ
zlX3mm5b4jCEP61BACj+BTbyiibqpJcKxVXCtLMMb8yxWwCll5c5Tz9JMlX9s9u8d9yiBxGgf6SE
mTERYII7PGy8Etd0Bs+YAHQVylYKEWe318mZ8SNJN9oXzAlcMv3jE7UC/p/SsRNllGkmRGoZ9iJA
6dp6HXcdB/vr6ImrRO8fehwO6z+kkXB5+Q48RRujNVydWVkfbT9XKRrgAiA8toPsQ875WtUxH/9E
zm2mPZRJsG+5pNIUrzHiA8VIPtQu7h8bnH7ZifPnij+zAT4ssnVcW5mYSeVDEWaYcxCd3pdrco0W
DBWrQdODeZ31xNLdsy3dFH4sOg65pZaOH1UJA1TJ+pjKcLRp3qlJEyxrYsiyFE440IQw5TGTJLHl
yDqfEQs//K4hi6Pzxe3rw5RY3MV2cHMJ/Qw+8XIU3CUR6Fwv+sIzzU+SmaHzeGbtsVTWSWD07hMI
38e8+t5wlFP6Rj92yWp/O0WhpF6eyGuwx6MJYRRt+Sv1RZXbiI73/IMr8R4Ohc5ycD+T0a35tPYD
wlHjF7zMX5Fgz+PPYz66Jk/nVJaRomM720T0XjHPBBT4DyiEoafgcgbxlrcsePjRHMbERXFDvdtd
y2d/aWEZPQv+FAAjr6z3i25mFByxCAXeLbOpyO+rqjL5hee4GgEJFRTsInGNRTspQeptJRjfCfEJ
9nAOcCHoJ41dpJ2ZkXkJgBmB2v1SEhqsqIvdJlBCqY4HURkQFyUX6zSrLOnQ2hBeUGbzwWYbGiU9
2oLk/l7Sfg3WAPeU9JkuBpJf1hhxq0cus/+xMP08igqUjW/UaSR3KU5dADDMuJkixozne9WaD40D
1PqBuB8N+K2XGYN2MrGLpKS3iUEKd7xXSn12dOzs9Y+Caob7DwpjmIcRQt7z7IyqkM1VHMxkToXT
1DXa4ru32cUAfbR1pTUBg3BJ7bPcezhiJfBtNvuNISsM6kCb0kJeRh1deI3LKyJ89d01P3ec7HSN
45m+V2v7ruGBBNYH+v2vpk2najJHZvh9eAsF3VsTZcH52HE9JiXL27j9911JWujIYhsSOrz45IUs
4N+lEeyf4RWoWwdXXMKQgT+CY/tyA/R7Rl0e/Wly/6e8RxxFhPdwC8pkeQZ/9eKIOUUA7aRXxiVd
4Upl+NpP0pA4fSL3Jplyf6mtgwY5pIUXLDoZcgRl9BUW/Hjlh+OPrK6t08kFcZ/oi0Wsp2m0QjRx
n3Y+XCIsEbYz6GJbZdb5aoDn+bMPQyu8L6dR8SBXJC+4gse65ienXBMC2PekEHUGgdobOZwOcLTA
Kzs7JmTIBITXXhNz3ohfWseC6zJieqI9QDDegyyDE5ars9JzR+wE5yBaVSpwCgI67jnXI/F4i4oz
GfKhihQJWrvySdiO3gt6ifLKF7FGI39KVlx2MgNYDMKg6S8cxKZAdhmqTErnqbveZak04DMijbWP
/SkJpPdko4dlBMhZ3fsgZw0JhJVsTUJrxKbsRQNtLv0XqwblvoqB8TmJq+ASsSpscAWwxcziZWo8
u2QzKB5fA/4BIHQnCXyB7+dJVdz/4wiIRsjd4GOKX5Ki1VxTGFt7U2qRNz2GgmCRrorgYkOjGmzj
W5vVuwNwKaLcxCEwiTisifrQ8IciF3SrWmLbErsYMdiFSywyI108kfUkPEyzRK8TjB7d9MyIHaN8
RKGYEpquSw80OuPkVZpb3vRqxoxZNW5OUxDDklZU+uQjGYUHxrrpmPdJVdZxL6Qrq5ylA/B3+R0g
vAf+gXqGvesk6/79pYI0fkwdRl+9vtyp5oZHXG7R0rTvvv/bFP5r0FXOP+rHSGQGwyISya22FT5V
byvnIUWhtBbnPe7DFtofpj1TDjuwke92nd/68i5zv+MEP8DVppCV2HtgJQj1Pza3D8gqPPJ9XAbu
0hcOf8jq7EmvmGj+LCeao6SPalampCOR3KkERwCmq8qFHYT8lM8bOXtjHiELaL9I7FELTv436JgN
lNT92B/iJslle6R4bZTGYCmTm52ODYsM6vn5KVqw7yhL5l+HyDfmEQSNzGXEcpkJQBLECr3NG/KY
lamJIEaHmQFIZq1VTiGEoaEeqkd1Fm0HIgkiJ5vS9md82Fr5fLUXAfB+B4QmpYSMbz9X2LOz/gLj
L4UCTCuPe3cXU9efJw4eVIeNkyITJVdqPjY2K0avbB6iPuesqL4FqoqElBLX4H/GIZBVyx/XPuQn
dtR8o21g/goyvgPVZlwfYErwDa3diVoOpElGkbZO9HIuf93Mxj5MDtNqzZJ6C9tsokNidZ3Kor/r
CE8wTpIt2+/kahWErRTiCc7V3mU0TFHyipINqwHtSsSFYXxsUHTRHxNPX/ISrpXoVBOb/207Xkvp
lW920JDx3SkyCogb4ghqtIktprCiGwqNw/JqIaDx2Z03e9ynQcF6HbuCTYNkMUWRB1Po7X5843sY
/L23oody4mdMeDyNFh/oXfUkniTwXohgb7hm4cwXbkrkDkoJqf7cy6ty9cU1MrGMHWqqBZkUGeh3
r3awIrvFQZlwaTT69LcZjW7ZeQcP/Z0Zv2QGleUi09y0OKKpLCZejDFcKlX7CcGAzyc6Y70TZycy
wKO+30vckmRbBzclPaOyDFi6AJ9ahF4bsHoEfoV1syrbbDyqGljcJp6PHkXoDCrRTWZhKmvyJaLp
/sipzG1SBYnFxTOa0mQnY3QPTGXzTecNlBpmg9OChhKYkT28Lit8Hvs3d3NCKdhIcojEjI2FBLCL
FsScuGIZPYDjecBwJlU/ZUGlV7/EJwEuDBJSpapQbBBCI5JUgva3mbh9jgepVYnLzPXycuJnTPIB
Ym/fzKLXrJz6nN+euXIgb5FygPnRaYzetx71R4ZjuIt5JcKQ/z/ipuOi8SS3raVjT6ilV1HbSXvk
GiQQKQPRQtsJOC8yn7dWH1js9l/pZLWMmbnqER7/FWPxe715GA8FXfhcdJnpckUdoQGBYP/QJhCV
EuAEI8TQSMbfJKbJbdQh0lTt9umrfbWysW7bfZq86xW/8AaRHcGwXRpynBDADhc3dpafmGcOUmN2
prb5xu6/eN/Om08mjXogB+DnhkyJBPOsliW6kN9a6TvL3Y8iodQsgYj+k7+TGBfMFMytlakSnyWB
twWZ6LGLY2Xej2AHjVnAO9UI0AclWU7qq5ni8kfaJqRqiJuE5WvF2DQdtXpOSGkyYgG3mBXNDRhn
GwvrQ8CWVeLqkxGFq4ZHuemG3hZauM7mAqM+vqjl8GwgKFNTippuMDXt6dhJR4MuBGM0DDOghpJa
N5/kYhprGJ8WmxtOhw7vAu/2+yPagH9k+JiBsnSkElOLyCc8ykqDnwnOiX8Ss9zZz8zQRpCVWRqo
TTUW0uQKThLCiiSKRPkaTKUSOqS5Fdh6OlS8974L7vMeJy1L0fNAugAVf6W+kMerpFGPcrUEATzl
B93CypJ0uhhGx+XLd881ns40C8iTA95L7kMPoHQjOPa+n8+uDqMHedyr0yG3DkqQXE+EhddBx53T
kCXiuabkjqJisEZcrvjAUgxBgljQeLZnwJAYsAMOCPCedmpHRh1pCbeDd9FUs/TMn+/3JLMEH+Kk
XJmZk42XN04IP+APCMRbZx4U+xmM9NYTzNK1TUlDdcp33zEwEoA4vh3KsoOP3NqgVXJXmFo8cTgZ
hAMB3p0DBMMK0pQmRsZxFt25zHAdIASic1PWeGxGrwpGvlBb3UJEJGxH6Ol5kUeCbkRS2lnz5rA9
fpyWmTryqFUId+AcG6Dj49TLVc/4X44n516H5vaV3PzzoP+phmc2cbToi5HlmjPiLfD5bslFIiOD
E+83vhN64JbqWEHuN4VV7onRxhJ/6+TA17QzT3qNbHd4lV1B2mS+DtT7MKKtyt3XWnFHU/g3ZFjz
JpaMZN+gvzCEY+hzzwQbmDAl3kWJipzXh7HZuYmc4v+z1lp4DO5w6dYgUNZ4zWWNhGpTLZaDPC/x
8/83L+mxSKCS6GGG0CfWa+gFXlMXQafIOtyHCkswESpMk3F5pkZUqxLldBU+WULAbpvNxH3K0GMO
RElpd/FDi+SIaXDFILKvst9B1vyZ4AdTQvAzO6SAMNqKUw5XLIWEdyAHKjxkp4pqU9/U3m/yu9T2
jcOQM1WmnMAZ+0xmoX+8Cv5HPWORfqpvC1cSM3MYIPlwShxVkwQ2k8MkazQ4SaaOMVEOvOyduqhl
Yco4tpr1WyceoYuAh1HzM2R7HrLIeJHetlQR45h8vx85ALkrh8A4wPHIJc0P7cMNJq1etJgjzqjN
Qoq/lsHNYARMBjf33R0y/NZODdMxJo7fkYNoMby6wKo54iAWpAQyLaXHyHtZLSEAMZVQGNtOQ+Ym
cPEqRg4RbDrcjJofUhfQNm/allCkZcQ/MP012jbWbWZoF5bRJSHUBh2Ik2gA4vEw2woA6I2mgJM8
pjj3sfisxC1H/3gKx4fFeIB6Nbu1bEZJGtI7nuQsiZe9vqikDwKS0f1Z9tXu7bRL4xEw1oaWwz5G
qY8xWb2jpJXjXC1pDLUK6LU84FWF3uRGnzXO1GWnluiAZlZ7R2YVu81d+AjGGOHeYIoIJbZYXyXz
vwUapVg+5i23e9SsMtRMaACoQzbw9xGl6/+U2sQ0JHeqwjkVb5y8gd+ajA360TOy+1Yxap8UpHSi
5/GjBUlM9wnjKt81mkIM287MNWZs/w/ob4EkL1RuKNpERe/QsfejH6gfltOWob8f0ZmMvZjp13Vr
Fzcn9OqXN8kSIpx0z/8qM0XzwWDKKlOESCiBDWZ3m8c/FDDLqkQpW9Ap047hgTs7bhsdK1Pz1cim
DmlJzoXVYpmlJOYBueCoViivOigh1bkgRjI8hixVM5hRu2NtBcblFlMvMERvjWqMml4Ogkiy//AA
MrH2a2WXMSr4nWcGop9nL1DnecDjOmohaqdWzPq3qh5znCOnZGouhn/8IFiMWbslx1ai1B2J3tLc
ByVuojSj//3WdL2cpwWPA3lulZagPBazvR1FsNZhKzuYnydBQ60+aa1LmFTVo6tmZzItkCVDrt4j
EgGx1Ra/jPTEaUs1t4mgSLbzyM118PDV0GkY/qxe36AYNxAflJGom0SNo1lgIvDNTTlhl9MEMLda
9ThdBK+3ru5aDp0Hacx2Hb90/Gi9LrliECczLbxrEmaukPT6ju2QSHACF0vqlsn0trUPwgQXHlxq
PaDKBoMij+fQNlCGZWHyKxW0WzwnPjZxgOAR4YfrXllCejkaA+cjF0QPtP/RmltCHQzRgo+x5Pq8
tWcZUigQ1oXrdHX6tZAwp7/RtA6PYZsH6VxHHDHBVTxLyZXrb2Q4t8fps4SBUN7XLTp7AoMR7d+5
V5mGLOetPYQPYupVrVJSSkJ9yaglfZGfgGtu8tdiaNs+v0gV41sLTEdOW2q0vVeTiJLtGvPRBZkf
hQb/FSIorWjpiANnyI29FbdKNbO9dIabOozE0COZkWwYDKkSjVbI5aJnUB7IBLsPHcKmm9g0NVJp
qXikvquxH7q0Qpwd5vKJAjAeCgBYH5a/0pA84gd/jtX8Sc9XENqLmzRWdq+LehF7ZkAglU+1hjQ+
B4j/sjBUO7yP6ziYiLluLa2D8SXILDnqHveh8VaOTzg5cPHzW9P7KN01ya9+Xbixi5oVqut4fot9
IYj42VXRtBq/9+Z8Xq7OC272a8i3j3ZBYMSS3XDJq60kcA6RBO3O4VqnFzrOXbScoYURU3yxFFuB
xZ2sb4kO9Xs561jvaJ6kLYPtzRAEfh9Eki3nBOtX14LSW4jdRN/ymiGt+y0/fKUuzQyD7Lv66fKk
CvzQhWkVJsic0Ut6Ntj2+71x4WgRFM0adqvOj3m4sf9vxBt5QQuGHt2LoFfT0KXLnmsBlrwvAdTR
m2YtpXexjCEomrLmqXuU7LmJ/C0lvXpvl8hYTM/B7s72hFslC7w0edvWZFFKhkzaFEiEIu6FCv1j
+nr4ZSXL9Z1BLuQIhmVXxA0zzkUC1ZGO0SEqL6NCS+OUEkH1bhAR78YE8H9rjXtg2RJgWWcHb09A
DiJeVVFLV1OTKyXlTkI0muKvJ6qpta+2vNWDrs+M3qVZMd+n1bgKG3THFmhzRnKXhAOL2nLucQL0
DIF0uT2yrK4uVVLR2u7C7HqMdLASxtfRPw4RrobIn2UC24yXRdBHwdGQ7bm0B/NQCYlelp/BnarA
MbuHTZ/Jpq520hmRcARqVUACsYByqEK5/4R7GsDLEjONqUGTc2/0b4RHbPpHfUyg11D8ARnNZScb
Zo1fZbU7HCb5ryj56AmO/fD3sghTfNfvKWTecScGFqVRkQX77mnR7uD4PsgxZ4gOtpG2JpNyWyOf
yX2H9Sc0Lt8llTPjiuGtjamZoHg22eweMwXYgYHXmKFCH7EQGPTCUkbwvgLHFjB9BI7b7z78bxYF
oYTJQo5Z1S9DYYCEQaIForAUW1zhw9Rx7D9ULFYEE0/mN/y92nsn6ZLPIU7x1yTTB/lPtALIZj7b
WKZhlc76gch54NfgBdsCJogwue7Ws4xVLZtLnpHgz2vtjwfT1lWkRyND85mAEwJOwlCLXsH7RtVr
jnNEekYGeQuE4bGNbZ7pQOz/kP8rLnNX7UXKmEuzHRhjyIU3m4w7klg4PtBsSNx64Bd6ad9jXYi2
ybs3P29zW6H/mx4oY97KfIeu1BvdQ8epMAhwxoAbjObK485uFyknuNBj3TyKbXw+JxoUEmHg7B62
4n4LDL1YNT1jHM+m3Huo/NE+/ORVvsNf8u67003eRsBdf/k6ZCfpJzZy2rSmJLrgmvK1ys6Zh0EN
UTH0oQUt2lcBGN9FbJVcn9Rxw6+ZSMczK+qRe65negP8mWzzaBm09HQT8Pyy0+szEwnoo93ft3qO
H/errFE+YRODFF84H/Y1sPsv3isFXFjl/Qu3F5TdBs9aFvTA0/PdUw+qzK9s8NtM6J97QAvkgYoI
VNxU45tctbE4gsCb5OXz5ji4VH2a4lQ7bGdj3U/a+ajN52H10/Z/U8LxFN2oONTwxU6lfucl6JqK
WLSXZQyJ5w59GmC67ygT4F7iMwzFLN5NqW6/XxNkpQGny3SEmdW7XH5UakWS27yVWz7OkjclFm37
6ZKS2iVD/9QlHXVEXzvIjZXlPN7rRDB07X5bO1xwRFUrKdqBcGfqu/PArRVNfo5kO26QCwiP3NsO
tr66EzAY7kVnIY+/jGKYuGlKWn9vaU+J9O2tXle2tVBn2BonMQvM1dbFm9mnuOd00UbNtBtpRph4
FPnBaBwShrcuOzTLKwTWXYc0jdEgJaWlorURod1THWmOtuuFXESypE0TZ+fapa2ar3Wg0GrSNm7E
SY/MSUPgTbeWsClvTBt8eVoDEkZTVoOjx/4BnbJa+FLvI5n3ny32h12Zf0Njk28897IOSXsHi6tS
0CbQfRWy/43g5aBFrFjR3sy5YhG0DhKpnLgR+YmMG7CAIWCU7BtQUCH0M4/QICph1oWzphCo0kSg
TDptY1mABBHbZBMqDAWsGFKC9B1wDcfeK4Z7EjTqzfJqtYYrDrAHT/ispMnTTueQT+QWTWAKN3Ev
zawvWyUzZY2S2Ap8bljOKFIuSkgY+oS9vW4K8h/cnu/+g3NDPqeatzapR686opYH2W1/xA4UMtUZ
9zHZtIjojWtOJQfpMbko5Y0K27WkyJ7vhA1LX2EyRIvK+BxVpVGeRRAzBYiKhbLLGbbqTo+kSQXf
AFMKO6pSVKznFpHzzV78xdS7cLnJ2QxAwCqsMDSiMT9N6jEFUamkU1v8MyZndVqInQmBThJODP+C
aw0txfSAi4qozWWQ9KDOqUF4K+afMjdrwRZg1oJptuKKB0Bg87Rwl7b2saxvmN+UyN8y4ZLLfJc8
mCsOD7BI1iit5zixeRAAxk+cJkFziNkxZX7bEQf3i6JAifbUqOqFtCdCNPHbOXV0VUSa3AoMjY/F
w5e88p7f+MiSocsi7ETww8vYL8NMXEfJO2J8Btoav/ILeIxNH7677n6VfcNzbM6apz4iTMnH3JhA
21V1yyEm4gc9+7CJDnCAkCaLo8EID0TmpHf3KvI1v11x6xDFPHf7gxgxAWlS7OPfFDl9kY35yDJh
6MQ4lfugyP/TgclAdI88HKfygz24dalOkxfdeBe2P4Pw1h20x5Ts6OrAlWm1VaZhIBKqPo7BTPqV
KJpwW8vFJL2L45FcmIVnvWDJV6PDAKOvt4dJAmzG4BeV8ErZo+2rM7Fx/F24DfkDKY/f4AYmaV6n
u4HMGiLVzzuLX7198Rk3q3BWo7yQ12QqeEX03WSOsyNZP3askWMbUmUzLdKo4MPk2WJgDNqc3mA5
duhsHMnJ6PNn3vXjlMFDEARxSo79WouxtCJIIUNpRq0RJ2BdR69VXfznV8bKi1HMjnSisS4n1ZYC
msmbX5guvNmZcyqDxsq+sgjsZkGg2CN2AyFvwE8dtaC/ZaDe0KYYJXPElygGj3mE8+gq+H+kG3ww
o8JohRc2TjMAmZS/dfewfpPoQtO2E90/GRlqfsfMxwvKDdT4CPlBbGjgdPH5R4hnyFRhRexXEE6W
+gOp64hJMHhf6hMKnxk7iqd/r8aguHkmgHFxIBx6sqE3qbN/Q3bYqdSKb2UwivquRRB6vSok58Et
2bTbuA/2wMbvj+JWZYlRR1wImXD9DQg/xh8wc+PeCWxNSqv65ov8ZdrwPq6lvNQOR65YVVDQkNFG
XS6072H8sapNoWziecAGCLHuGoVaoBXd+DREcYaKZMuNDqL+ENmcJ0LRmzEq0QSG2+jmc7HykdSI
4hYwcYGlutjuiOFO12yd/61xXakOOVj9GX57cM1wpQoiX9eDvxhTsEbBK6ycnKMcbhTJgt4jxc0S
2q44whNeAAdn4wSAGA0iDn44LZf/wXoPBkUHugqxItT7dqZD2sCcRM0Ro7xMICYC6drtFi947Pb1
sHKSl0io3K9nIGpMtUX8kAnRPScK2c9fDZJH+saaliH1Nde2IYj4qsPf3bHxqB0vhEWvHW9+cCnF
70exYKk5ZxRyjjtItFtLkVcLRm5FSrpIuTsa/+4X7tHgInuO0zcWihAx5bz5mBCgTB9b8hQV/Mgp
7PsBDsdmYuvKtZJD1IZII/sGf7DgYEBx/Fpzm8+ZamCLNxZKMfPVe7BQT7mFVxmPa6ZOSQ7J0GKt
q72iMWld1bOikaWmYV5ajwTTXI4Me4NcKBBrSHDvrip0PTdxLhxqYK71jqCbV3t+CdRZqeeJtZNT
RqpkQ5oUKGkKdLuV53q5kvzy4uwOHgoPBABW6bKZMbdDs3MzypiDgoBQ7MFQIN+WxIXy3ZRQB2B5
4o/BurXh4QL98YYAdBg91buHbgztMsfsGtczll79L68N1ETwgSpMCpgjOhvDLrGMfSdZ7kULdLJx
d6XyUhQLeqeTAL7BWbpqD/8fEfyJxkC1Xyz3Qx/gqeF0qbhsotu5caam2SRRPwUeq4LtAhYjBOlj
l7VcP7dARSnHEST5ZfKMGeTbD36Xh4CVWhpdXhnZjBuvmQMqqpGy5AmkcFMpGOAwPoxOHeeBh6kR
qp4sov9h/6oP4o8VbgR34aZwAQoYu+McKALwSeSt+QkRHaeWW6WcV7xnutbjeHvKytqoC4lfhypa
RBcjZdHsn2YntRMbeHd6Kuuw5JP+lo1c6Xu1fXF7pOyQQ6qJzHTwBXB2Lt/zmcaM8CfIwK76cgYI
7bY2I1wWk09TFpK3lGvyEPFlGSc0YMJ62i/nbVDEj05YO///PF7agOeM/PkGk0aj6aWyo1YhIgQC
BDpZdVda1KMaWic60+BqC1cucHzguiX5S8VKTGUIP5zOnk8A4PqPHeeMiyRXf4SFAzAq2nG+3VDe
NYQea8XRaLQd6HGoebwCepWJaKgTL9uIcMgW3oXMLLZgPm5BLY5vdHFgDpG57G+HiKKJY1JLszvz
h8iYUC86a7WelbfhZdE8+oYT+lfEKj6O3jotdid1ND2cQYBW9KNITT71oOCYF8PwQIMl+6jVKyKT
FriTpic9Y7jBq1B6IQZlmGAv2NOrWnVsfEtH2KOZBLoyqG6KS01Zn+XoV4U2lGIh/piSPcyRe+Sw
5cqs1j7NTy/yyg5ELJVRe47yX21ZIS2jiDhZ+cLXNntwpU65ZtnFPJbhKg6Q82lUoJDXSbSIgDVS
2A4wCwfIz6moOtCOhJ2hgnmkVNw7D4SJp2eACIZU44cNwlu03W5E7yuwUWZPVpL+6qjNU7h62hkR
6/Zwcdho/LPVH8lGFP3g7Es83URtMkA6pHMj3lFU6EfC4dDJMIlVDCxygzifGPM0YMCVOjtPaHU2
f0g6OFQNhyH8PNXnkx/FiANinViF1a0zNnfZKDAOc0SZvrvyEVx+Bs1wUUutuSkTRANU0JEkWwEW
Q/Bey9b3fLv5AX7+cyu4wXYKwnAhjB3tkCCMtKYCCizTaG207NpeugtiWg5vAwaXMHEv2/LkB+U/
3PSzzFwfcxHAwUVT4qLRqJ3vQHfu4hmb1FZZdW5S6GAniT0Oj4jSHXQpXtvlh4DAyJ9iJ+RM/zYB
YjwoI6w/Ou/dyp3/GVRp/QAWxwPhX68vXKNNoD0rOMcpe0/bgKXay+xwS4rbKPKUho98CJsVqmYH
WCgdp9Hbx4Audqu6kAVMSgG0mCXWvh2gOdZJVCpvjJLe11JnhjnLQ6xkHgGIAav/T6ZVXSlVVbqa
RHUrRNNm9kS+5W9B+Ac5cbUDkoM1zBsZ1HMZmAMslEXq9k12bQKow5net8lrVdRRqbBr2keOJM6i
Ri3fvfHS8JgHJXUOANnQVZuG6jTg5rVqAHxjDyZVH8XWC1CsT52GvoDTaQh6Fx0nnMcrUBZ7TNt/
B/2rtrX00SMVUtg+feDfblyMpeplBq/kWRPqrAWhcaJyyBgAiLsvLC5/QzEWqWGiz9U25T7he9lE
FRgli2+iKEetiHz0ZzoHpiWrHPv5/vSSDkQ9SeWicRGfxFTmlBPqqt7jNcPW82BevhcxpcnDfAJq
nBXhT2aX8uaNtO9kaQyPqMN+wIyEmycQfNQzh6peqqEl4gUb2SgnofmCfvge25T9pDztOznUwias
aXhIT/VjHw4JD3VNOVvp5lyWcVNjj3fFeZQkVJLzb2ikcmObGOAiIHld/iDjSdKwjVZj3AOy1SGX
XRGhg6QyAwpAy3cPZK0gx0FTr9C4UvPAM3K6gOJomUh8CmqQHgctc6uh9ga4qNL+PAYiInYRGyWM
UgeQsLzqNt9h3QFf/1fA++idQX4uEc3USJMvp8HeXEf/9kaovMIabpb73kNa9SfHbQvQ0sgW6Hro
Nh/dw3gM5yc174zSn1ldT0VOTFy52IrhpsnoH/d/AcflsanqybpTy5heLTLl3Vsjf0+f/YHJdAYQ
oPrODS1OO1SPVBp83J2j3WPh2+EKCYmGtCg+FOVgy+BGvGgxPDSpWIsbJjlUrCHAytwRBnUCqtl6
F2flHRR6VMWMfsB+l9fhklFqqPWTL358AapBPpOUdyd3ky80IjrnbiYv/NdpwqoUUaPPE5Vsa6Qz
bNdIfd916xWjmCUf4RbwQdIE3ME6TgaLr597HoGsjZGsJgEQFEzFOQD6p0ntvxUHe+rWlUN5UyhX
uQ2OAj4h0U1MI37wQzj1UYU3pApVnLhM76SsyGhkSctOT4dcjxikwlYOwgkvnhIMr/Z0jLgOmnWm
21qbBRLm/xowqF3rl/Vt/YUF8XLo8VXw6pznDNelAAZs1jNkJfZPM0Uye0wSqh5QxyWV9qbW2xCQ
x5mVjbwWmEg9WkVLp9+vDvZYzlK/CqsEVb/un0JSh32LAM+HaMtgbZilI3muiWHBY1zuY7XcfOjg
gMxQakFzJ8D28kpI/4Xba9/anc7GaTyfqPlny6EiT8Gru4+D05rDGjKxx2fMYhagKIFfYHtbBtdB
Qx4twDcJ78eRpvM6p3bybemTtWDNKm6xf65hWzcWH0dMCIg7mN/KJUn63BHXQbq27qOdkA6Mb7Ks
p+jP/N8X0xolsRtLTlV8QGMx0Kpo/CX2/LwHOCXe470e/3cOX3i036ipZfDrMZxRZ2VH+uk7eand
OKIAI6ttqcVDDHk2MKSoAteAdWgK+qjEY5EXtqtq6S69v9JuzTwvaU0ocvYgC+eDU6MDWCqy+MwI
gHn0aspNR3jgnT224a8Vs1Llt6a/fp1jTblVcTpiFzSp4xRSyXKfHvvMB0Hc2/LiDv8ToiUW9GXY
OAcDI02zAzDYeHCuOz5Zg2TEsGDXTUnIABiWRTfnlbW2wRjYyTzaiE+U65atzjXR4ob/dUkdnrr+
S0wPLABscKTzpvIkPMzwQT6vmPPxkDs2eTLYCVG4I3cnARdhQMIwPHV0gDIS73b1n/ny7tk7LnC5
5SCC8lim42XyMEb4Hg97ogcorw0tB1OFpzylAHllxYXuCLI/jrdv6k9/AhZAWGRGpKEaP8wIbdo9
txPX5LzbamDchxP6HEU0M7AxbLCugWvrrHbdxJXXw5OxdvqTMfOelPZh51+CldT5ILcUo8W7QCRi
6Gl+a66lw4+AQ207Id45pbzJTiPgSxaa8z3Bme0LTL9AyL8LjGyDMfGNuDtepEtay2MbHUA6ahQE
GwBLRUXjyjoGKb2bIAkVa1FkOLOGzPkqjLwYrsL0vz6WIGsgBRgH+FT94x6/wTFStjRUHe0CeC8j
x61HAUL5xG28ORnuMCUFKtSq6L17GhSamXWd3x5thMwT3NdvQF2b5eVmaVOuCJcreKQPYqXzo1Ut
GUhNCn4lFUFAWaM/zSwYzdDkdX1C0A9zWS7t9LEkT/sYnkUiJLjsuk2TTI2x9OAoHSYhxqbc0V5l
wqkIUAou2eiEoRWNgwvMgrkAVwJY6+/C4nDNBtRXSYLjatHpjwJb9ZUsJdQXsQF+O3M/5uOVeqEL
LuAXLAW9/fMZ27t10HDuCNa3E4OCJ2i9+EgWztmswLp7wZAPQmQsPPoEL6XN36Ghr+nOR9ZUmynl
G7poSL/pSAWM9PRN+NsMdDeBGZ7UTBWXYtc87cmPcxMQLhh7bnWmJoN9O2N4OYd5y98vFCqONyXC
dSqS2HlMOYsAfWIuU6qMxLIxtnAFLiYqqBFlz/yHyDN0Zw9hsR2T5riFExuGdVUPgpPEc1aDElOG
M6T71pYpHkOq1HM4nhYpNATO+Wf0DdUz10R2i7zCTGoFfX+vE1/Erwt+Xkbk+aMVStEhzVlhaNv6
4fZ3jy1DQiNsuWXO104nPtLXVt97/p1Ea2NjjsIxp1IGcyY310lG8UlBkVfvBD/mvjQKjAtMp/rN
W9BgiFsxXl/eA3fvDrCHUAZLjZ30ni38zjWwvRy1NMAWLy6Jl7wFMLndJjhb50A8bu71AMPq4f1F
Kunmf1b6vmvZrksHeWIPMXAYUryLo3ttmoHfjcYcWnvUyGOlqEVdZHqZpkU3HCK7OUOMSdmnHopN
gx/wIRMZMqBsBUvHEr32a/4hZ6k6rVkwfDKYlwuFjLfp3zJipUYJqzllb+vAQjkxZMA2kIf4kYM8
l1HGm9vZ2rCliK4pG8DPQKxLnH0E43l0Kbo1BVsZzm2iYBYRBJ1udyeT3vJJixsBAAiZndCM8CO9
11VKv8I9ouhfWwXlAvCsgkJd95C5BbAk0DxXfP+3IVufRZXzJeE6YmGI+U5xBMQouFTrgilCNk5p
wYgvZ7W/A98k794MA6pAiO91SlqUUaJKdE8utq+hP9fvOBkj7q5qYFfDK9KnrzR3yoVFzqm/QjT4
hGca+kF8UB2wmMHhmbddK9jnCET3M33XTI0Ic96lj61O2dN/dbQmarNLMLUcbboMPE5Y8RPkqg6Q
HsUHncyE6JQ3/gehY1gD8F1a5E0olOJ0Qi835WyLvrthx0c3nqOGMcQbvi1Ex+xOFeHnHx+NCiDh
LMedEQRFfR2aS7sUsgmhq22KnJLbx92QZbLzHK8lsKUxhuC/GcgzOCOnE2FTz9NXWKzdPYwgSJI7
jaRQVpDfhXrsPnkAgWLJiuVEG4yHXx4K/9WF3mJM4Aj/JQOMK2F+4XDwWPiWoptOCOxfh88Xr8nK
Q9gRdqAes4hmerIOnPRb/8h1Y4GNBwNwHLkH2viL5uFozNRr1tme2BvoaTfPh+gaBIboX/WGBYlT
LRXWAHKcy+ff82ffVrxQUF6MTUYUupAubfcMswiVVTZNs3m+fNkDk+FAnynx7qt6RcNPGO/nIatt
ds3/8yBcim7CiZhHQDIn0shNddNXTPbsrPmh/wklF0PHRo6BBAKuj/x3I+8KkOjMQhBDjze+SGie
1fEA3fAFwrhT6DQ1Y5vBtMHU1epc+SgQvg1xfqdrG5BYfoYpqYritMsAmKEbsDRNaj1/xU+ef1g0
dNO6bImFjePSoyn6BTw/KUoKx/OkgR2UXvBdfe4yQVaboTftyD9tvFjAI+iG5c7XroFOpcf+ml6X
j/B8EuSBlLs5OL7NESZ/qabCeJeWuAKPcgo+16lAVdae4jvoYxEbB/ppfH8pXhcqf1Ej9xTKei2K
PvDm2TTri8hlMcEDdFjkIpnWdz1esZ9XOfMo39WEvzKkrNym3F+5Rz6cLCgci0/vKimrMnk2WMYK
mgbarlglCLWXw/dDWgJVmhr5vfjdYF+f9SRcFMIfNEtkTp7im/ybkIdFpfRxTp5O8/ydvidNzPvR
tk0ozc64iJ8roEbY0cvWAb+92cs0r55Sxb3FLgXVzeatkpwL19B5hoV0nJO6c61mSLQG4kVohzdj
KL+tJVZVZ++as3TZnsciLoiLHIEgw8VhB8EzAvlY/cZAcw4/Izj9dYa+1zNFj5hYp0OYf5eWOG+m
0g8Z/XY1KGMubQ9zBmjjCh7TghuPuXNhQUX/yXhZbtRvkjkSjUcrEOFW/U6rTOeN2Vn8BoTcZwAK
2NNHhoMPPy3bxrwvl5cI8wZGY1y4XKUFXuWlMlrjnYoidqUsoOFvKst/Oee/UpjY8WWFY+9KfkrC
nKUx2u0ASIcGQrtcyXHbc4UMEJGgLugQ35LpCEzf0HeQnS61WvyUDvL94IwQkUG2CARPWUaG+jlt
z/kQP/1QfJAydMTKeSx8hwY5iOMhDgg3kkFEdVKwJQ1VcF8wqijUw8rNPGtRfFTGrp0iAmjrhBW4
5hdlJCUmmQANIPLUwb8epj4Wv5v/0g4jmxE7pI5wYCQ/b29CTDEGFq3+SPL/8W8CEeSrdah7JnyJ
BY9HrD11LB3XO/99WOyXosZlZyhQcYJU2H/1UA+772Q1gHceSq4Sho6mGNkHbtu88ewn5QBLuBpF
ahjNwo7f9LuWurZqIZShiDzD9zNyqIDBbm9bWURoC9cMdZhrP5KoiqfeVr79dqGV4bgUjTEUFWX2
zc2JatlQbUgwgRZR9xZHXX6thDsB2WJ2KaxZvLk+tBABKxyXMGsxGfiUE3+MlcuhIgLC6CP99pTj
Il1OJFF4pTcMTgxLHMQbyUIJpbRjJzjPKNBRruc7fzdAoGhtyVb5w0DYF4co+cu3UmRcoD0b1nz6
pmQ63t4q5P5gG61+8ZvF8Ylyfe0djTsS9eEDjhhv1Qd/wvs01Z+OkrwVCda0/D5gXmpFkvmsM1i4
czMVW12p6NBXHcmR0CKF28w4g/KxN6yi8KNQU6z6HOWBDljlE3Ko2aApYLPKAm2G6Mvy/O3c0RBU
OD34BXXsIfTnaKqWOGZFzLxgI+Jpw34DLi7skR4jxxrTCc2/xqAYBWWGcEXACRbI7NjWJdVnq4bt
Q9ldBaeW22ry/WQRyutkaPUVZalksJJmgcC0WucxtsRI1e1O/DbHcEQMIGnuHVsrhnpWFrMoqRn2
srE5dLL3VxcYIeqOy7O+k1i25YmBD8C9UbNTMg/z7HaxYaB4p//R6vVEn7Nnh0opxizh+KjueFOJ
jXU34kLpxMP5j7buWjpt/pzve00Hjn0q3qXFnfvqBNe8Jj6EguL81RderT7RMF7XTAIQ+HcLtacC
rfivkmC/GcoShf/qX5E0KNwoJ506EK1S7Bfn4y36BKTetXiA01oi+EIFWUrYyx7m920MwKbAjm3H
fIi+Rk7GRg5n57sOAqLTloT0Up2ZFuTq82APWN64CQvpoT8iIxDOzjycb4zTpz8O/N9YrgkUCjeE
H+wGUyBY+vs+F6QcnGltMYuZYBt+WbfkXTh20Z516gAJ2W91r7m5lbnnc/QUX2CzIPx9T4IxsOU9
8b772vZsVvExnTMU48GNdfMR9GxLDCRwL8H8bgdTYxzOakOeYnYJDEpjXd/aE0rubEJMWmVzFjP1
obMeKT0KZgKQng8GuMaFakDN9dOGryCT+2P1d2O1WYep6vwamY2rnqkPqW1g2KtY+CF3WUJyajNS
pT4WD1VIAC8FWzxTiqDe1mpilE7NZoNFBj3OpL6BycvQjszwIGHvXq9jQ7ydg9WHoqgsa6ZGa0Bb
etOGfXfshsFg6yNVfyjgFQBuHq1996oDVWctfnrUhL0mykJN2TbXF9OlGt5OfNe6vhFybVWwN07i
k50To5GnIgOMXlva2TK/BOkouZic0gCAFkdqUfzAsVO3FqMz3SKgx9+wJ+UxYfeWeOj5pCkwZTKj
o4CRnIlG7cOgcPzKr2N3ajLYq87W1hi3lnEG/c0f+35rbVCjz9fpYGIarUfvJfcy1zFpkiqALZwn
MNz3e0RZaXkqeoRPySSxjM0+g0FscgGitInik1gpbsIjGjjrrtNWNX7mYo7AdI4eZXNeYSneCxs9
DKQips/3ui1Naf53IKgFhrzlsnJdwiNpdprhSvcFqIgrnfEXvD+/4t0Zk0v5Ru06+PafpJqEjQmE
n8foiNud9H/XIrWBau+t6SjrFyDP5mC8p6BUbYtoKZGrY0KVmsxClJwwKc4T79Z2yKHMi/dk7p/S
tgtFQ4WQE7Qsw9+3CiT4fkvIw7grd8IJsaOc19AM+XPQK+3poB2UF7760XMXZMiQf+pYlkm+ynrW
jHT58VmbX2LtxMZUbbKc+ivzP7JD+ZLJf/VZr8/QIW7+zuXwuRuWfzEstcnaf9hUzVVgykTdZR1A
Yya78qtMs6vmNAMeAIhD7MRwC6vZwhrNmBQeAQ1G7wnze7qcgkvJvDysMzg1x6R+yl4J/BO+MlvG
LRHFu5YVP6tD8ZtCbmeKaUaBYcOa88ItZAjEHSS4Nqw74CCmYn98WdyarCUzPCCWlOIT+CGhgBxE
lzgJ+nDXcRF0N/PhF805MD/iR8LgQ2x+fpXsxVkTKy8LkKEIHIpJ6UEPM1x3Ei1ZN2jLaKOY+VWg
V60Xy2up3bwAOmW9sWA+5q5Spgh9d+ko0Q+9XgTt4oxbgQCsjFkTr6v/+WVO9W4cPcvWfaiY1fAe
N2KDg4o1Afpb0qa+nosA9UxUpHD68UfWCspUOf6i+da6zzQ0riUFSQ5sYZC+Xmu3qu8/8fLkvIx8
mYlx448DGMZsivRshYHaC571iA0i3VNWwcFcv50HAtlSsOhYIYgF79JDQDb5K4oS2UrHpIP1Fkvc
Nd6lN41FP++lWlYLp5qXnKeGNcm0PN7TUB5TC3rP6phQz3Z/CVBhQIG7EY4fRtDBK8t337KgQ/C+
eRMNrM4l9ZD30yBg5/19eFmJsBRHXh6wtCe75JVr9r1Nmqr+GUU0FQBTiJw3Yrbpctb56LwN3fzW
ApIjrHj4s9y8rAZWLdG3ataMSlKoFyR7Ihp/DZ1NuxjbZWLInkXPRmcRp/BLUhdji+ZvpAMAoQXj
B245sEbwoZrouHjiLBqWKC2IB5RzJnh7pES2V2CaqTYTP4N4Qjk7aJJsiNo8a7Bz2OH1jhNjG1BW
e+1b1mZNaWcED+MhmIibogb37FdhGCAxM1QqRrjt0AeIlzj+ueNbvJYquRPTQOdizjNioHgxwmbZ
9w+gYSu2Iob66n6skFpb30cXZmM2qpMbcg38Bo1aYUj3tG8u03QHtF7YlX9b5GM+CRLg2HKKAPyn
X1OL6IAdC9oztLzOmTmjWfvbIn0dJlE+KliKRpY8NiPAsJeVXWsUmimUryfj5pkO02/pkHAhY7Q8
oBk9hFUl/Awr0QMagb+b4rowAY2gRbLv7yqPY6C9QkmulGfaKGzPpZOprgm41cNSlkDa1SCKqK28
sfAp0NqHHYe2OHUmoRBfD8au0bqOqKUOb8BfRdws2nOpD0wlsdmM8PuV0u8jVTUqYDtuWalfvHzU
NnWbeRSdkm83iSg0BUYVqlLijmNJ3OD9paqcXb4608loD8eq9DmfNSj+a1oP+qlBRI6L5B3XqFpE
Obqc2xxHcZHBoP5lMRC92n/JRs95Yw8oxTZnPx7A9tuAvltL9ZrVQOGbc9Qgi2PwDQjzhe6h7mzF
zi2SwtxgGG3AU7MYaY2kA+ShtZyutkfgSSKpuoTWJeWuQxQGxJm8+brpycTDWKMlTJrF9h2oh31Z
/5NydpB5o1lXdNBrZWSaJVSp0xYiWzXeGdPQoUesSxj1+L+72ZGp6+HLmssjdfqIsd2OyafR/3kh
7CLWtCbJfy+yBigDrJEvH67eYvZr0XihSDCL8QYM+OCOZJIJgQVJ255YYOqzfxsVdl4kTFuhO6ib
LeeBJ1YvR+M2p3w7fNbbydrJiipk76dtB6Bo6fs9AMZs56Zq+i+UcPJfXmD9g4RIC5Hm4u5go3eE
o6Ve7YvP+Se5s6fHDyMITled9xfq3PXLsXHhzrSiwBDrVrFUDeUchnUPn2SB4NCzRJT5QAsJIzP9
+GLidU/jE9XB/CZv7ETtAb8cvob7cpBligNJstgRaQn75XS0n3uLGCy02etU4FMmOApjyg7Mpnd5
RX42O+OYZk0DHQgmIri55oIXVr28JukDPgumypim9bH2iSVV5Zy8otLM+GW0lj7ZwN57UgOevQnj
8vdOboXbKT4HSWNWBOVyAMlxdoa+Pe1AmysYdEXDzUFV5tBdXEm7HKDSIm2Zcxihv5YADQgC81rn
HMOvfhqzgFOJnOMhHnP7p8R4oXg8FuuMPHzZuses1NtQdbBVPASDBvoJfc3O5rxDlPpzJj7UYWi8
+we1nLDbzY/dxk61/KcRhIX7PBDP8wDLfpoO8ycKLH4MF2602qD+BVvL4xFK6Ar5wYyoVfOegxLV
GmparfNnRKtNj/APF2vZmqR1POUAjh9oq/Wv8a1zDUM2xMoxDw8II7/6sDzCl/iW01Ts1HyDW6fS
3+3w2YEjc2+DZvXCYIINwSaZckIdVMKnBJhKyXhwTlmSDREmDbihMbZ3JdFLlHTUu3jXFTEv2J93
GcCoRj5MbjPPX4gNtPlIXcE2Qv5YCOqRum11Q1hYqORVPmIt96wW9blPgQ/Hcn3g0MrVQ+a1Bg+w
1qo0c60IZmRsG/qnFs1Tk73pq1mbzDGzOaqjYAmPDzhO1ENbZkaZ+OiNu4ECXiSYYODp+4AP9lgF
r/uFQdar1jajBhp/o1T5gy6rLT0Xqdz8jpULgL1R+uylgpHAW+lrU/WgbORiwq64tvDYjyZpTkNv
fLA7iEVxOcU1bV0dkz7UKOwQ5pUeXKNffpu9Qr13B9u5CAt1PjIhNenxYLxeCSSYrxYWhYvsWJgv
9ngUWmWV9XxwQtaq835FjZoRIw9IVcFZB+u5pFJtWZ62Ufr8UdkNLhtjdQHHrSZd4U6qOBYMMPVD
aIRo3WHNUE0ikV6A9xhs8oxw7Csq81laSA3MGcr+jbveysu+YuCItx+pOeahIJMRrlE8yqmRbGmj
Icb2lot0G4z2leBU+dh5GqBFvPw9hhgis5FqBX02P7oIrSB9sRSsngrTrbS3SyUQnALXtxceFt7l
fCB58Xv+oBOGGH4nQSuQnfwOL9OzqNN+Nk38KmwT0Ecp4yBqfWFxBA389EB59uaUdiopSGMHjL7/
MOxugy3CDjYvI9e7iQDIMjdOjnXe6guOq5EzUXA4oLvfi42LbHvNpoGZofZdOGjDafKIUTf27Rga
jfMFcvaAqPZDl27YHxE1Tqrim05EyNqIJ0Uo6e7kFxzMnyqxOQCZR8B8ctdvkYxXtezy1WggHPbd
ZdaSXTt5c4YuZU/cdcsCohWe7ORfn9JYtSawbhkER9od25deH5tZsajc56HVxBupf6vBo9ckE82o
BRUb29P0az+Yu0/bOq25fnbqtEwPh0OyGO5Oi31CZOddauVz/4pEmyGee3Hy5ZCvTGK3jIB/Jx3t
SZAiEWCg3rrjJwFBAtiY4jYq33suFDSf7JAaBH9pyYkQH4kEsCHTtx+ocoe8pZyltJn5e4uGrsnp
60IHb/vvblOvUP4ZXRJCGj1M9Pd98iQb/55bnHl0BYDJVwZeChTFfeg4i5XV2nBAa69Ta1AJmFkF
2TgTEZhyAr5oeUgigxfGgMcLhDWeB4i9fURDeuiCjUuCY1YJi58eRLtidoRw5UKlbFqymmnUs6Ch
dLWOgHRpvnJfP6OWCqD9KtkLygKaecih8UcNXOT6Nib05v6tPP6qGmna/fIHo1uRRzArf12XUOeG
yBVV09YbheY/oWPEiyBbw/tlgKokBqgPaset6vn4OdbCBAk5/eKdJY0WBktKfZG9BwfOTa/d8Vjr
dT3nlUNf2hf/o/gBFqfKOkgZ9p+OpkBCJ4YaeQ/t8pN/6/M1E0kQAk5mkSWsbdSPa/0GvoH8maOh
uFKYZsWbTt2AF/TwWBC+8fkMY2xQmB5zyHWrqu5XWtMj3z5qinp0CWm0ZiQbFhaxmqC6m19DjgvT
5/CGbHKaxBAeZRrySV73wgZZUP6LN9O70tchZA086NifBo8FDoy5MEkQuHozXsD/gYz6QRiR9jfB
RL8HymEGa6p2/vuRULQaJmHi8s7wV/Tfcfkpgd4dCyDkOD8LIOeXLmI1pCtnA8zBtl4fGnGMbMG5
sZSLx9qIxzwsRc8HEBL9CkznkA7Avl+26V/TiOoHyITq1Lz9NvSPmvGrhdzP/YW3oBpIVybuTNmt
8+I34JKZTVm3OtCYjDNGkgjnyYF2SvhACmbOdJA0s7NkTL/c5lExnDhVSVoGUzUlK755Eka5Q8FQ
lzqo8YgV4w2Q4ogGYOAusY9X1EWMmjktPKPjRP4R5Xp6kWuencuDjjgsQdBVELMpTO2/6Cs//uvf
r7klrUvFTVTy6/Ov330JPR90IhBOClN/GNkUqFSVei5xAEAMos/yJhHTYv/Dd/rSAoi2QMb3KL+v
0vP8sUVz3aozlwbPMdOyk48yOi/NvB698d3aznQZ5LfnUM8I6QcxxTuCR+k2P/eMKlP5vxzb7uUa
tpIBS/jszOlcOpdGcSZOAVwOGdNx5Dfh1JFzSoGTv5Ngs4d6T7C0FYEu5UtwYwgl4qWL5YwnvSde
pu/RGnRL0sKqF0DB+ZMGlWM/ducagVnX1/sCmeEMAximxsKG/X+EufjOW2OWWHYmw0a02rAGNOkk
8rZ2ieivf+HPmyUCn6N6c8NCSTKPtGpV8K0WnSNGrD3OFossA1B4+UhE6SxoDD42myZY8VAgcYQi
qYcuM6GKwExLZ+llunLDXvm/24fySoqQmgpK+9BAmNGMlNuHsggGq0QiBnu2ydYOIlIVU8BBVG4b
kXFwlxC5SFKOK5kRcToq7bw4lkWfCzLPlbMJOogsdaIG8nrKBylM4aCOYHxVXBrpLPsQn7e9U5aM
lsyE7P3YNypqFOEsuyd6MA7vBPI5lc5li4rsdlxLDTSn6i92SUYbV8xC6Dy3hLm0tEBoI1gK8Avm
RSMuZ9VFhwmEr45IWTTmlbiGph+5A6eXaS5IY40MnxNkyzVa/2JQJ0eYuppSWKQ0iO+voG+Aqc/t
gqc2rnSBUbmH4L9gbKE3tMG8jE7uWmmRp09sPWmO9dRGniBxo9rTiihDG2N/AW87WjT8X3Gmc2vt
5PoBUs8ljjCtDTDtrx2XGVNK9E/MI0mBFLZ2dcOx1PMOO0bGXZx8yI69ueCh6So3WFC327ydB9vT
wuzXS6WKhL8axVJXcGnfT09f1f3DFeGL6uTmiyhwI4rMAR69QqZa2p5GJXrDYHlZk6UOp1TiQaBe
JIEHMT2zB2UMFZwzpGWR37cIMLD5hK7zPyVOQnP9OZF2fnEy9KmpQ/vAFcKPzVKpumukcDtPMMl/
qC7V+0SnSNFNpVHTkJkYcbnZuUmTNi2qb+jfzVViuEF2rGihqRclalNSNfljsiLRZHmVVolTzc8D
BG4M+DpZRHgIwOdGc51PfQIqp4M9uhvEO4GHFc+NBHvJnDxWPMx0KIf486RgFqzdPkXdSqeeAJEr
aiY83O9mSrVp1P9deE1Qbnv3wXqLfCNGS9OLn8dNB9zVeipFMuVQy+0y83ecX020SCjCrv5mCsu4
Z8OPaTPxE2ZoQOmdjB25VXHjsXwXBZHxmO/LlFjHwnnfRoNGBaBs3x26fs9NOy5Eyjq3CI5bgllz
4bYjT1i4JLzhs/OP7J8rpYudrJX3cnVRY0RV6n25IdEBUBdlPR9CuR+/BkaqQI5LWQRx1mTupUu6
WuW9zWio944s4b8CCK7xkqYmj1a1tPFyC57XToiauYugI3tjT0obImj6LElZkW1UF8o6SJG1YBvs
3jKXvBAyHWiH2Ak8EqtKF16ceygLA1/3WGDIGx6yp4TZuTNbgwWBmJ2PE38haC3RfpV92RMqMpx+
1TkrdnhZJVAN4d5iew/mBgrWlPIW+ZSiaDfb2V3/GYIrB7bkp2zeZgKX8lAjz7rTvGP+zDXAUKay
fRLweRyqnKb0r7+DuRnqL0YYF5S2fP5mLbsGVF2Zqxfql3/kMW/Y6pEQqUepn7EQSp0PYQRICCl1
T/LPdXe6We9ME8GRS3SuoLsg387elrjsJiEHHE8II2ifuzP/PGQotMDGCgCN75K1UQdrsWT76sGo
JNkvH3P0CZUco9snBOaNLVmdphlYdVZB6MNyD71oJMAnACahzogGVlUaRTC1+0LXyn1lZPfckJB0
jHy4Xgata2QVF4cQ0+PVLlJtc7njLpLEfzG5h+cpIi6JpXaMUmTj1G7py90BcaLx6CRzGFGtQq6S
P70/+Rk8KemckEY3vQKR1fZ1mqdCPOepdSuR8uvaq2NeDk+NGdh9e71ksHsohy84Bubm43al3CGO
LKFLg1dJ3y2j+4gAVNiqgvynpItZjRstKHyp0KG6+dSpfglTzn39iAVAJgzImm8P/5v3qpReFRMb
rSLg1XIstcpsxMBaGhNSvc7XHOWZqXUTTmwRyVX/GickrlYBzT4Py1R8tumQ1Xax9amv9J4sp20U
f13vRneY7HJNb40EXE9mwnCPvJtsn0vBX4j0s1nswoJNpPedZAUeZnGNSa1mbE9cSxCTX8PG0gi4
QqmUchWb/IKOwQKU92kIzAtm59dWBjQdxDnP9r1uP16+yr+KBetFjR3wRAY1I5BlMnO8PjFNEahw
c/479JRLastwFKKqtl/eO913PMiWryKYtfoS8TEW8iH134WISaz/uh9Pwyuz/ooPmdmOxN9NvTs3
wQ5EKwP5L68TCHSr/ouddZ6mtP8NVPHCs8F/hMMkzSW77hdm8x4MLzWiLOIL15Ux1lF/vEHEbAyT
z96OXLt2ZIj/a50lXWOKJ7ZGtJGm86Sbv9Eo79cChGixjaESAfuVMDhzbcfGdDPOrLpBBtBfguEM
eeLaP6LXwq+jXrYNtdRe6Dp5RrnhgLDtUdfoo9kwVoNkvDl1R1o9kE/5xrdidKLGP/r3V4Hxt/P6
Y/e2GuzrhgltdK2zXeg2OAQy9FFXrzVPTWmygsIFAAdWzOBBIm5I+1yRzbR8PrfZJx63EaWefgZO
HDG2aDkPf4tq4IaA2Nf2nrssbWB4GpeFe9jz4XqQeFRxVt12Kqlob11e7u0epa/vPNb2/R7MqADa
8eDep5X1rWzlzP3BKbU5d8NrFxgSpYOf0jkG6KJAxSrnWOeua284AWu9yWtVFHOBPHfg8GP6hpyM
R8J0P7qRJqkOgzhBjjZ1U1XnwX9J3Eq81DcvMRaNnxmgY6ECM7cS8YkFxnltY+R0TLtEdKhyBFm1
s9W5ishUv/9G8OfDbOcd4iQCRwJkxNcHGt1UeIhJbgha2cCS2alBbqsO9RWVmMh6qAUrZalyDvPK
Qe3ZGel+vcw+rozfbfvwoI0vnw2900t1viF8fjqSTKVPsCjDARH0u6ngQ8Tb9D0FccqsEwUOrBn/
hiZwzUKF67dVsFgJJdmb4UH9KLs0zZaftccHMwuAuPitGCLzK2vvysX/H0Q8DPP/xiZBMoUxRLcp
Zx4GOJRU5yAybj4bR8kz9wZBc/ph16L2iM7avCsalCZZGFo1LPOUBKvmZDiU62vz4NsGwrNNSwUG
6v5GoRjk0kf7OzDEinz5wCTHYWFgQQ2bX9QMYmV/VKelTvLfl6DFmklfEoDoPgQIFalPevzPreyp
r82KGP75dpr0hohNIBxL0ER39X9wi9DSPgyEf900CHmXpo8q0g+RdSmPnteiNUDm9tCaMNNroWkj
knine9a4Jdpo0S2Mq3kkOM3sZXpP1JJqli3AI8BB/Asz0UCRLGsn7wLAyy1KXW5oT+tpE0FWKdhI
CuKAttZrIhSqsG2hjRMWrqQRFSCyZs9PMJ2oW6jtHWfh4TojTWGvvtAWY282NX8b/qXFFIK59Itk
4a/Fyno+HliR5bacGzAJhg98qapYE2Q15sf9NQOGNuv+qtGQrm9H6Oq4NmYABfHLiAbUxXAeU+O4
ddD3LnS/E1ITKsEnoCnD84/4gLfuyLF6Wa+02a6fhfVYUxpP17hibP5gTyzU5Ldlm3mnsWuYpgZG
BOY4iNEGJ8+xtX71oRnfGTdW3Voi3F6zdwa6nJb0yZgukhgafSRlsjIgCFAxASUMT2xxmWCLLbmg
4FWRG/Hm3XihSOaDqQv2cgtMlifxF9AK+Oglqej03rr84l9qIPFdlFvacsub2PwnIgvBmB0yYkdr
ON2DCCPY+p4TBOFLFBTvgL+oth15b42VPJhRYzcYuaSYdO4Y6mRuHfcqK+96AVVzhieldDgBzi0Z
n1OKJtfcdcjD+wp/XhFC9rl6hB1TACeXUyfWjNt2u8E66yU7CepqWI1yTyo7De2MQeEqsswg/F5G
HQuZXmTpY2NANsdZm15LdaWd8Y3mcSbjpfD6fBkk76ZuZSQBxnCE5GRqzVABzKbMQGUw2vUeSYJV
rdCQzzybI+c65kRUowX51Mh1x5P4YiPTI+nLgVjPAoLVtHy2IxJ+RMiT0tG1nr3dn5DS8C3XWCs4
/U7phyi4HstPM7r08nKIs+HJY/y9/i+7i7SfHSfJVfH2wn+fFjQ50diEe1xrbG7kh2inIXjsVMbr
6zGu64wk5P5GJ9okBBDlJVGb034c+w0q/SlRSk8NKLdgZ+VVz1wh1/B0yG8rKywH1/OMhGSUMqBu
2urHvu3Fdb1chIQhXoGkx33mGgAEreGu16MSKuGvJ2IdPmGr0/tex4iuqqlaroIEPe2Ps7NUxWa+
dm95GscraoJk/ez7JfjwwEUKAu/CKYiicd213zhcMY8CkyG1KgWRfacOdlPueKf1S2vZoirbVbe3
SvVHfheiicAZYWUFkMSOq/vhbabUUWTRSrdXLfQlX3iInHOtIeKp9wgjMmjshxXTWUbm9Hgpnjfl
Kzhyxwd4rLoR+eT1PbdV0gSOR6u+zjNPi7yG08fQYLw9Ag8xF2M4yPIkhqrcG7rPsq/GSocJF2jV
NRBrA+wPgOdft48OyBcQfb9nIPzrbHekd/7VbvF0NBesynDMfyIo6eByMJSbfZFHheMiHnOYzjlo
Y83KsQYQUSabJROVNEkcA2nQKC8V/Bnh8AmcX9pR3FD5tv6cUtIbqCdyocX6fmk65rZgn7d7Iy3e
5yqrjp4zbDKsoYpaDmjNRIquevHl6/uvHtIamdxO31IlqWgtB6MtFXTNj9NzYd37j7sG04Xq8G/r
Ww4imKop4B8GlLgjbm31ZHwr/762UEy91eRoS81VSE3i8Rj578X6bDw3SSIYNEMZDu0KF63z7MOJ
xBvGjAXZOyOWeqrHoESo29nKQ+1ROuN8fjwJ6AvmEf1Sb6DrpGcmSA/0EZ6TMOSDUwYGT2TA1Uw0
Qm0o9HDTwVPXUNKtM5Lm/mpRbW2hMpH0kqIh8XpjPUXSeISnexkO3dAl9NRkDhDuqieBuBL108bm
x/xnSdVefxiCl3iKSkr1GJgdgYLUrIDqnp/IBuFTe9p/lfoJO+j2VbdUOqt0OexRkjAUeQkzuuqr
ZGVyDlJ4zKK0LB/brAc+HYnv6PNO5MdVBcdWpO2UxoPJVn/X1k5DQ6YfA3kw3WYSQ3iOrlg5cBk3
71n4aZIrYJlzQDSNw+wdWW5sbC/a/GUfjM+XqyvHEFWdfVlcY4uzJbV6cOoO9vN6FBn8S40Y0zfb
CBSb8y3jPdaGJ9FamlifZSfHLmCQlfL3L3KJfvqB58K0CxCfX/cS8mYSI9LF5ZdahDX7y3uq5OzW
FHcLtmiDh/CDXPTwrhrFIPNQUgy3DCbc2Ucfn1glPlWL0B6CARZcTp4AFBzpjd0P6qIcqZQebB6T
uH27AD54CaOpknCmvJvFuP0SlIrOdARb9mZb3TzYqYkwVIEUTqcgVKV8GFf+LyExY4BDBngjRYJo
NJbdy6V5M8Ec5wt1cBufJpYwlTSD5jQirE4/SSAtaZ2xZYQO9Mx9AOfoBC0fyaeaO/4eHaVk2GFY
DnE17EJYUlWFjHn1hsmrAaIINSw1+m1zcOzKGvwrFISmbhTh3VN5kMuK86Ns26JQBJT18gZ8ImTq
W08bHlUDVU/nFMsiy50/Iy3vSKYQonFbiH/+yjNoHh1TtVHHU+6IXtO9zLATV2qJjveTAIZCNTQQ
QU87T8jPsn7gKm57CR3X9QNfwXZyFhZJS9ug5qXzqjOtiTd2NwgFVEgbjryAy6YIiEbCdvvelfk5
h9yVndgNDENqb+mM/J00OOHdpdFWwc6+9daYuV14s52HYjgPVKZrxS4JJD6YNpU11n3Rqg2+9AGc
aaSbv5mpzMB94SM251pf6se9J/RVJAym/R447h9cUFEcWnlSrGzO2l5kDNLGkEFjAAQAPSAeejsa
8mzSoWYo1oi2wWh94h8QqYVeS2PzaeWXd6WtE2xNVNxOO9JU4esAgOYYp0uWNobZoyIENSGmcNLW
O55+JPFkVeTo0bRakKdlUUEQjBNVqedJCtwFI8M3l8NnXrLRMkEXFMcv5EHXLQwcgGLN5lqqj0QT
XfAjzrWt1LJqhBsoDsHaD4yJE+q9jjVN0wg0Qox2apsA6mDklJyfDOT2b5ifpyI5F8Spf6Tx4+Lb
zTrbH7Y7LjQ/e+ZE1GqrblA/xqkYimGU7RTjCrxQXCc7PWeH8jIMVt1EUNaMT8qFxtcuSRCnVmBf
OC5LsIoKYDQdGHOSuIU0KcEgPNFKTtMZ439O+f+TD4Vh3qofcBUHZSmS4MORXRjBiSOTXv6M+FJz
xxWYrMzKGO0j+Mh0lh1bqtZAAmzekgP+RZ/Atj3oSxdX0iuHDtdUT/vG8/wur1257R2Z1QkbktV1
VU+737UIrAR+H7EcI1TYhdLp8tZHaSqt3XuM+pQt30S5m+KcO77rpdBOLP80z4h80CDAhCCQ95Wa
GvH/mJjaoPPy1DRKQJlNi4V2vVIulVeDndRkdeaSCmBaY1Ut2LrzFEqmCtlZLyQg0q6QXuM0StTF
79C+vg4ib9J4ruXkHNXrW0Xbj6n0Lw4WT1/50BheLwM6nfeSF4Qv4eaxZNdIn+Fv0/QEoQkvFpBf
mFW/k+F2ZFJYNfRIogt3zWVfZtWE8z8te2ByMUyrW1O+fcelLIwaiyoaxrMxEUQ1chMupzsgRrMp
AJDemSAuZgD7wNvoC1AJU2RS3kj4S+l/cLU84uw08Jk7CAHKUkc4wUbVdWqb2WruOHQNxanu1SDH
hZflZOXuh7pN+JEQGjPWryic1yKVQBuxvZdfg7aVDD0WSGPHJIbFDo3Wsj7sqCeCadUuuTYwwjzu
Y/VJ6kRKibFQIxXLbeHjaq41tUVzEP7OR6w/rQQoaG2tdXZ64h8mgMLZ4R2SKv0fSCvmUCh5VzNK
nCJYEa4blvYq6ibvLZBauCLO5CPOSKNVsDnlWLmY0KgzN0W9PP42XPqOZFI0v9Qc60ADvvEpRBMy
zAaE39QhQobHthmysVN4vqm8GD+INgFwWE62KpxI/M1MfDWy277VWxRrpX0MgEd42V5nHFGdoJp5
hYiNnbijLyVkSBy8FwoZpcm8Smnx/G2daysIDx1PB1JPyc68CjNVwk6Oaea768MXTIoXOS0nnPhk
VOuUbrWG6paPstJ4aqi7QlvGUWbuLkoM5uVGuMwfrnQSeRcf+WmL4NJuvjIIPO1NbZyND2Qt0QRe
vYWZWMuDHYSm64OvDBgd2bq2S1oI03Z2mHyO/F5OvYgTQ08XZGxnpivUPJ75+O49gSfaE01TBJef
gVs5Y2GR9WG20RdYLUnFvy99c969unepcQ7+MbbyJy48maOj0dCybx0WcAYr6rkhv9dwuD/SGnLj
J5z5Mtq0n3s3/J5fBwDOQgu6ZcENHk9hzmzyAf/s1/IPnuKxbMDP+I7iBpBCa2BDtKem9rwc0/K5
COidizWo14Ji35Wc307hn+9E5el08bObeyq5bWbngb1PBw56lVKRKpaNNiwZN+jDKcQ9bgiQ03oF
uT/y3p9RvwncFGw1LSZnLmjm/yOkKSkWhc0ExZbHv5sNipgfs5s/FOdJcjMsRsVxm/piioTAI87W
KFuhVUYzZxNkNUSzXwPw6QPqwITw1g8svegmUj+qkAM8G49IHHnY8UAf58QyOdz8z8N9Vo0I+CbG
J9jf7YTW0Be9MSEIrjt8mlsAjorICjJL70LFCVB/b/aBtDJJBN4RZVQRrfOVBhwCBYkl7JZuRcEc
Xnff0Fjsl0eFbHOHe7/PMDD8AjjCERGVEOY81krrPHeAyMhpAZVc6kkPf6kpFpzvVf+18s2LicdF
IIvdIHmZjhN7rq8I5xICHfp0+fP4aCPC1vOJbL5+3OJAXvrXs1wy9Biaw8A+pQhc65O8jwsROH58
v+OUZZzBRLtEdEA7khfKwufj7c+kLycAmc0zPW/EpO/dXdqm8pyMuLMDDb/0IMTZr8ku/wg/HobK
hayJi773KPyiba00akt5zRiKBQ2go8gStYlSLT9yXbP+lCTKmSaviquugC+QY0OXPvKUJyPBeVWV
tyFk9ANg+Z7akscPkdDA3+CYvkMlUaiaCSk8CVWBaeKuF3vz3DNLt0BT4wzIxnmpFekpPWenlBol
56wE2HRdwtbNFZ3RQIZwveBs/fMWUBXi/Pgye8Ia7DRiSU/vIyXt2Twvt65aCWskG1SJAJJDwGOJ
Es6vrJkoWvZsQrJoAY7Q+tJ8EcV0t5U7gqfmiQx8H7CORbApbsIImUSijKCYbaWclJQOJ9G0x8XB
ZrgHdwk3KFvWx8Vf7TOYbNit02YEC1kovGX3/Clw9hUXYtoGALcUwgGjrI1SXCdyPZNi9IsFudbI
Z/tGXRK/LbE7vJmFRZf1eZkOrGmDCZhW/d+Jhi1X0fTUyheDxNKteE1zYI+oNKLxJOnqK+D8ZJiX
HOxqtTgYw1bXKSoCilblI4D49+Bfr35Y/SF4V+sB6LXl8qH2kAsDmCinqVWrkr8C4PXxaQoEv9ue
jP8fMZ3W7PG9+aAXoeHAttitRXOJSU8zYtSDeQPA1rWdd0Hf2yLb66Ui5jQubz4iwtxZP4w04tBX
F7O7zi0qtT7S8QWvu2++IxL+dk/oSxE0cHjXOvjPdLiHCigHZVh6HjybC9SLAEzHPEi/foidMlvm
iQHbCRbuSM0NieYJqdp8njDjgEYS4UJBRvN6aSt4w8c+GbGauVbCdAxSkeyF6I+qO/41ZQUSIn+J
B9i04rSTJJMOGLoc+sa2o/cK/q9bFAQ2MpnAYHG9Hox23/DgXSiyfTdxeRN7kiIVLncYvTC0jS1o
fLL+rBWqT+4pln0v4/NJjRVLfQ4obf6rIJEa40hajJynSWjbzeu3x7OIXr7V8bXbsSUn6RWxtPzW
9upQ651WCMNaOIs8bIxBhzb2wQ9St2IkaLLniZWF/mXROHZgjOeuKi5K8KOG/7vSrLRE5Hp3iZKK
U98GUvcYOEOZUEleQO/23wIm8WrraRN40GYV2FLleR+ckLl2bWERKIF47aetu5iUrFzcp2MBYZCG
m5/gU4G5db1eE55ai38j/rph3U4LqVGwUZ92VGCCe/a7UFSQe+0w2DwW0BkI7ZU0CL9fOOwsQxz8
ReSVyeiE5uebWbtXwOewLnb0ykG/hdI+wehh4v5UZlYTlRNNy/nXJuK9nxtAhzbK9hv7ud6Y4V8O
4HDSCRf/7AIc7eIGHgz1Spn7STR5Pby8C1neYlu/ul8xgF+xZfgtq7C7I3M2ccwryQXbkPTIdtIS
F8nL6Aey8E7v6Jbl+jktxZlssQKZ6LfgqTwE6M+qfReoCCU+q69C3YDS+sLe5E2JlTqFlyW1QgmO
rvagCRHfBuhE5Vlmpo99cQ8c3CG66KiC7qq7LrCKnlmuOTOJuO46CDgPfOcmfsGt9VNRsxrAohSZ
wpVdbkVYbZNuN2Wxp6WS7+OWPs0WeqGrF/XJ0Y0fe9DyQd4tuo5YQ9v4eMbOgFDEZgg3E9vV590G
X7LgaVCZ7N63OpV0jbx3X5CQb8n6UOCTqmKfKMAlT0EkTgHGN/krLPdT1J+c/FFW8r+zabhiQk1s
C5f7TFZdGjcELQCa1vOCHPZ7C6LfPyZnC4zp9Qqux1NSFTEIzBSzP7C+oNwctJ5+8QJPgnRCHXgG
yoUApvvAPyfuHASbpcDEehxkyKsCJN7AbaesxJnFsQn0+eGZ3k0KZE8AIITImgM96RqAPsHbxhED
TvpIUZbxxCsmFTLNrH6VY8jZWlNfOtBeEGxHF6AM8tu61hAFZJoKu0VwR0CUPBXI0IFCq9u/uRFe
2u4UV3pnuDHhCkduRl8HpJ157/9VgX7PPlnt8CJMLCmYyJdGFAGn/Nq2HKNvEKer44wBN2adzYud
U2n8vG7cloZEvYj5ttDKKeurfbZZKmOgqr80DqCz123vDV4//67cPj9xQuYt5hhbUcJRvWIOleFx
jwy24O9DPNc/zlvPZQpF8rbW1jGCuAR0l6MKt8ash+t2pRbzCvaODwURaBzGye8icNJwwLrPLEe6
a4jo6j5vEYijUTxL6CSEQD7fxmzvV3kzJjDq+ygEFrydjkMenJQLRfW4OnkgIDEx6+GopbJMGDjS
lYM8GzUkfDkTdbhPaPWG76Ns0aWKSH2tWjm0rLVisQnKW9H8bT2XTrlFq78Yt7mlmulkeI9PXCWI
ZNiVjxbcWxvDOvGiZI5F8R7Z04eHtY6FLxHDvFM7fnZylyqiJoTY1jAjA9CqyeYoLxXFBYeXiznq
77UmSONSxSZJbZ8VqE6UxKfIEWtgJcqzjZkHFr3LWjbjgBz3DyukVhVUeJ7nITHUbQIH0WlsP7mt
4WCverzYSuWOWaiz370xlZWbzCVrHDNWlqpqfLL1shoyGZ+kOxKMZod0D+BxY0fpTixsacfrENTW
j6UImHlPapaGPT7149Gz/luzfq3gaJg6HPNCHrQqcu1E76lnTv5XWDmUv/A6AmvDxs8KLq3vd1E0
fuaq2flCKV2rQ/eeAma+pTgsiwx5B/UKyau7VjoDEHs2Lhh5HFq2drE32zEwkn7J6nN/SJqo3wZV
Ft+EXNEciYqFQBsnm0gM4FSJAQqzb47ZmUhkp3uQ2Xb6thCYobhCZ6WM79wReRYNNEnGUPn/PdKo
ZAHQqqht/QkvqlJTVbc2njG5CLc1dmjfj+KMu7eJr5AYiv5oUzlEghy6ZAJxIruEkbvFCsg6Fx+M
7auHKcnyiv1+8y7jGiwn9qt4FYL5Lk11W8slrVQfoOU8y7oXFw5iRiCRTxrgVuxHxJmNFuN39nyG
lunrcsSiNKmCDTgV2Tz4QPjl54Iga/B5yMvjbXJsG4MNhGPtyedzajWi3+9TQx2qO9eKrqFBIPH0
bK/ai3+e46qXwaSo3liveYnKjZU9tqcghyr76N3vu9S6W6ifyoA0+BAzfDYsqTEsI8rnYPOHt18O
S0fEOuvMm7t8opx+3UzMy7aeO774eVNxAsnVJnygb8vnyhvI5kr1dG9Y8cjp+AyhrZuqipl1VuiY
uZZ8c1hXgGI4jwxFTF4v24frngueS9nRULJDWnWlnlAncuZi78/84Q9CFi08kft9fFCxiX7DZXCO
zWfcGlq+ebsuN85okPmkVgei/0tWeQQVmekxxI333MseJMqqe3fPMqNNjnwvdfbiaHpy1U+FsvXw
FkKiwKxtqfvoTvF3buJneiEoBuxEtBMWTNx/HILW9GVEs1AhTl4x6ICZMTtIBL0zgoTHbryNBh81
MXLRNDex5QGXHpCKL3Ao6OwjSxkE28rIjVZ/hIwirP3Lnbtoo5bu7eXqL6qILC/m20KnGl5OoMIK
BU9x1rCShCwL5o3qcTwzixBVu3b2kCkltNJYThXRyHLbhEvuJBP2udKSv5U/he6g3fwHz2kYDugT
x7fnwf1tPXwjJCi4WJzuoaKXr7dEvmnwLU9HhRstedZPOOFdYyO8b0Z4EI6xbxSzPeI4xzCVe0BO
Mqz2g/d/BmDxNsK7Qc3YQEI9XyKHzEhL7PsjQWmh9kZkmVo8P2q9eRdSB8tBpAFN1bgqb3jlCyb5
Co05DBOkr3f2DnXr8Qgy2No6SRIghybPOw5pPKuIa1HZgaSpjff5GXtDIsM+MbKG01L4Yi6KhrjF
hM+qL1SApneCrZNSJ3HqRd/iEjh1+gU6VdvBTpB+R9l8R9R3U+S8y0yPgW73cZpZjnqcWkoij5gC
RGDBuerW9FDs1n4U90bBVUREi+yydczqta9nV9VqPd7j9yk2QZzayHF4FGBU+IyXwRxHXcucMKfu
o1jvHZAeuQeilk/RObrbg4yrjSzbhhDQhHeZlPz1EzgPRPzk2s3AzdYWE2h0nhrqGaDdKfAso3s8
7AFbz4ZoPZ1dmGWcZECrbq3bEa/h1ERq07czes5NHhdQQHMVZaqBYN4o8Fsm3+gSW5UjrAzIAbLi
a2UDbdAXdEofeDfju0+P1pzyUr1Kxb2xinZg9ZVoaSq1bUSX/ncSZe3UI0lyxMXdd+4evCfjbsVd
lkKiWIuE5tH/j19FK6tsO9IcYQpo0wAR/95At8ws67SRQUenAk60tcPhom0GCit6lacf6pTRT8yx
6boLE+IRKUFSUXo6BSLT1tmo5hirZFzYx+J/2OjTLh00RN0+qDfbGVDHabDPPqFvego70tafAJN+
PY/9QgkRwyDggczd6FNjWZib1aifc6GdywYU/Vj6OZTeC1K7xWptAEXAputY2TNsU8+NFX/wiN1E
TWEThOxcrhVsnXnXmDNmVxnuuUUAaotu1GksilGyAZbSZS4RkS7QLU48CgrmwT2s5vER8VvkjpC4
UULC8t5kkGSZPAfxbW5QACSZqNfa+Bakn1tEsv9gpyK+sn7Mt50ZfcaKWC4cfx81DBjge7kUUBEb
x9vCMKt8gYtFz67PKTdMVOreNVnCiAct9OQPGMoG7s2uPwq2/Ve/804q5uxiLRr0WRtESOUCIWrL
HvC8uQ0MjqEdvQPymBK5W/9gL/xqg0/Z7mIh26HPm0jGbfU63vyXXO7gF8Qvkr+BgHVWrAfH4LI5
Y9EpAImRjXGRqeqN52qDcWjsSdi6nO6mN3bTKywDk86PRst+VokLnVcX6cGdNBxGhujV6rJqUpOL
Jt9jlCY5nPCQKHQLN8diJQGoyxKvbPkM4uqRS3Rf8jcdmlVamzPr5Yv0rXr++Hps/5bfvKGw02yc
/+NOYmOYWDtwUS6CjBcV8XuWu0dYg/4omDlB0An54EVZu7Zn3U456NIZ2WSoi5cyhoIdMdLdfXNN
cnH0lrSnn2CyGtZot6CwF7WOluU9tpBMd+vZMA7q9AUmXadbu+fND9P+DEMiJENGSUtUcsKdBU2E
3SmkfLsGShe3waFDJOolh2Y9RsNfqY/oIWmeMtVzJccbn95L1J1kx6Q5LzMF6dlYrs2uxTzsvClR
IuNkqqyJwQBp/LFTPfjZ13GcalTilltpZ6blBjgrDYlAjv+0eaq+YK5HBK+g6wUmAlRK1Pbn5gHR
JJPv6wOdJZZCfnDZShaRcnuqfdeTcvY4v/nQh7ajg9MHV2X8aAE6zVRlO23uXw+mhoFZhdv82aii
PMqq6ddEHH55Ej071zLZVoVUjvQhwKYfFyQNql+Z0jkYA1HHir0Mm5U3cHbXB1Q63sy0F6e0tpSx
pqIEJltIfRmrDc/krI7LJN+SC8ShR6/fnc5wON754FJerPpU7pSst8Okfr6NU5ltabKT4rDNWcJI
9A8Ik9MWRPfevU2RHVEX2kk5qtvKmidHaaExi5N2Muml/rKJM/8oxzCMgNj0mHHG2k80BRtwf55p
OKhxn8bg/MyJUrw0B9vqQu8V2rrEAT5uqjlgVWHd8YI99AKSQrQGKld2wtVQZI5Hf43jyYOQXS5m
6NMlQeGhb9/bpVdkJg3tIJZlo08zDd0f0I84DIdhh4hs2mElB1yP8ElrPtg+/DDIhAsYiQlbvHVq
QLfX6xJL86fsBS1agF3n2RyyZu1i/utjzeTafVcDGaN0RJwbUSUGv2R/7Kl266cJwdWpN+OrDFLU
JbuYMawts4nJS0TaLs/A6vZS8ANG2SWm7o27OIIUxMAWkSak29/iHjlgCNNLbEma5z5cJ3emD94G
vMicdBztfxoAOWaoKC+mAsCH6ZrdnN3YRJ7eytorPo506kBNgVX3se/7NX/61Yjhum2fNOaiIBA0
bcvUwvWRuADTew2UYdd+4LzNpKz9t3ynS1If8KxTQK41dRtPMBj5SYj4LC4/eoN+wQCzSiUHHq12
t16vqlp+SYxwSI50/awk6dpx/hDZk/3kand0v7zUMPxGB6Pqh1iUR9q9WYyuaL9Bj+Tn6Wa2yXq4
/vxOyCpSm15SM30qJd5jA3XjUaMYfWKBJZ1LHV2sm6YAT5YBGItWm8ow3U/lr0JqoNt6coI09B6Z
3fFib9SrCh8lq846jUWxJkn9iwYTScjk18mT84rjECix0cnMZel+8WoZZzyO7dYeMRPh4hNZ6Ym3
m9ZI8A1spB9hr86HTiGT3CMrk+Q5YqzMD0t4+91TJvwkyytKL/REO1cURBUaD90kq3RhkdcVKUWf
HFTEGYgcAUsCHYohQoLbfTeRFFTop0AUJkjMyI9GZRWhqDyOcmqVs5LhVG1/KIQJC0J6brUWHN3v
Bs9AEWbrbMMgCouMttpTzuPkl6Uc7KjrEDU5msxWnS3tKU+emQbbVCxz8NTrbJK9unJuwqNehAHP
81CQSRHIqHQRVU56BkTswR9L00I1PzVpczxza+w63X0aoFpE8XjN9aFrPdtweO/j9QvNr62j5PoI
g7PwZvoSsvxJT2Oj5n0b0erqBFMBYQzw9qbp1KEIqDIysaGN497pIP7A6NBhgG0YFrYwWY1Uz/WP
rxKa9HumrjBeGmRIf28GHhy7eXeR9Zldi7+FxLjq07SFwIPihd8BM78eYwFQuRF5ePjvQGKci3zR
y3rJlww1fFthWIB7JLc9BlWz8bllBWbuezR+0BilvqLiSdB2sDAEVNW51zJWQQQQfaTvwKvYY6+b
FLIiDSe0/LSsu34imgc21zkj+vDT8Hr1+Hi/nk2eBGgdzm6X/JIBIAMOpWu42pPK4XoHNy42w248
CXfqUi0JTXD7/BPLrfUJOHG7W+F/ue+S0/zm7M+GLXILNQsGSKNPgdwuxBKVHBcfDMjgeqQ/QvNv
9AF0FhnLXQwaAtf562wJa9vWKn3RYZMVpKIGMn/0+0h4VSD73sfGVZBzxKyJnM9KxTuys9wUme18
N/gc3Hu9FqdHUQFn1GH6oFL9V3OdECh+3Gg6JlWqrkmXglqdmzGe4bdZ+/frkLhejQPJS7iwYXGw
q08FdYT/UEcgHDnQZHARKcIS1IyjO+MzF4NwyzPYAE8rKmuiX0IWQnrcusRJd7c+2IWwlOdzEFTW
QF3FsAN0v+VIj8PC43lw0rIrTGLfsx4PiKT5y29UbJO/fIkS7WisVKZEH/LjyQ1VrAL3zi2EFEVW
j5YFZ+rklU/X642vXr+hO8JR8ZsokMjSRidk0QtggLbyxEZWhnbz6jv0uMGchcRJJfdb0qwS2kM+
6BU5U/Iu/C/Q0nzQgPdGwH4YTdY5c26bjCekUO9H/4rf1iS2EVhPBmxPDnZaz1ey8an304nCQdC4
zWlt2tCC34CTDIhNdMQWjD8Sp/2hNxmbwXe7VHtP6blEmBu2GMyJslkgtM2nYKTyfTgKTXJYRot0
aOdviS3qdGlQeNWE9qMTkow5EyRVgpYQFZiUiWD4II0hwyTKV7g34Rlm241oBRR1jyBnhPaopBfV
wxhXVTQrI8Vgjtxc3aKBe3UO5SSzsCMVg3DcWA6bl/GGBcSDy7dBko5hsr30Zn5OEOJip0bwIGg2
2Z93f3UoDz5qn1MnulpryPyGV9noLnxP52FoHtczD379p/CyRbxfffw47VeDmvYPi6Jy8QAPNtkN
3PswoeXvQX6Uwb+OhOq3CIpfhAQxAIqVV3srA8UpNY5V7Z2GGgrJkuIwFo/jM6tDikUoRyO4AkCZ
Qt04k6um0F0L//xp8XVFc8hLvJnsondcCRhl6KBkNi9JoeWIXN7pEngjwy8RTDIFYiY5M2L9Z1PT
0WLG5p6i9ItMKl3j1LAp15j9J7946wuiJ8vQfTzzrnIY9tO0hm2HqSC8YXBIKhMkNTGqzroZYXn9
sRi8tkDx/R1N1wQFDwjFrsDMfP7DAsZYCRxCR2yz3QhLI+WkBiCvI04pnncKfdQHOEEKAETpJtKS
yTkB1rkLaWDVlDH06Dv6AbrM9EmS6dPchjO64eylSBn07HLuXEfdb50SPTsqqt3POoAgzrxkcL5C
issdk4E72Oul9j9hg759RFBSoobGzeakM3Q8cOCHkRsGIpyGGagr2cNSHXMN08cIiIsDPFhcy6uh
cods9r5jU//ki2rzABCcGClLDROuWp340kmbp2jFgU1zum3NyBx0CCj9nWz/5bDYxLeDUrqlw5aX
MN/NQ7hag7weU56b7Z9iUo4OkVwBdgoS2iGTggK8gyxAfrmN92kIgcCSmdUFzQpH0HbbQkgjJG7s
ombcCQrpf01VekeQ0qWxKONSuDtRqfMV/UmSN0L3dNBoISD4iQRN40Sd76Sz+lxKWhbL4EA3/N/F
LBSjDdrC3D8lYIl0+BS45E2Enl+SL/t4ApxQKYK6TxgMXtC1FEU/X5aav9ErOT262wUrPtCBqTpJ
a8p9MolQmF5EledRFpx+EAL0T6gzm6pBLL2saVx/+1rU1TqVdcGnPYINm2frg9jRra7zAy7jRxqs
tNIe0pT4eX+Ky5cuoe/mGu36rXTvVlMwvhrTMlooJgUtKowjCvIAnTQZ3guG/GrnlFjlovtVDrpC
Mf43j1388RoF1O5AWvVBXBJS5XeEgICGCUS2eaMwzN7UU4oqEMdihwgop7216yU4aLDpgzeI+ppd
HWoA0tNmcDXwaj64XvS7A3o6YHvqDjSZ2mTImKe0lGS5NjaJu8sDJG4SZ+B+JVP4maw6vreR1qUM
WP73vyEllaKXYF17BnacjtWo8Yf0CU+Yg63bqIhAPLBK0KCRmzzWQf7nuuEnDX2jTmCREqvFbtxi
FWY1kTXivXGv7HqV2qnP5/ZktRebF+gCD3wO07spr9QLP+WkpDVMZYDvWYCJnk3/Jt8AZ+UD9kBc
agmezB2phfpjTV8/k6SHH3hS0NXVBzChLnPFSn+Yh2Pszw3wXhekLrAULcOtEVKfBmCNtCieQC8M
2CI04Ok5kQWTxaZYmw2lLdBm3R5aPtabnGupyyQw1cboUW1UAJQ3ZJ6c3LoKFVGLvGMqbBi68fdW
wa2qvIpaEgcBOTpoGDfwb6QOLu4KGGsJhCDJnf22371aV2Z+dwXRoqNXqvzHnDLYQcuWpW3Cdyja
j5IXbZpJS0IIk5x5zF9LKDY36RTaElClNb86/mr1dToD1BKMEBPZDI/woZBhl/WkrpA+iaY4sRSc
xgejS5GLXmpJyvBfYp5ojW2aWTHCVaP+K5JjKxCwQaCG88jBIqqqZGI8BzGa8FEGaii1nU3wSR52
6QAPSSReEYMoQ9fDTHy2G6ZtPe1wttSxkrLfCMKT/Xq+N4Cn663AgGUzRIdQOj0sCEBxdiq/rube
Q2rzYSQl+xZ9R9B8K5KJU9pLKgP0lqKnCzsb50w42e/B2QNR9H92HZIUBMlYbozSDhldyGN8QUQn
VcUOqkfpUS6DS3CHovzZVpdSRw1JE1rGOzWIV5xaLtDwphh0IhjeYm472ZD5tS91UOXL7hvA1/Ev
IYtF2arZCHWGoTJn+ONfXDFEfmmTYhMCs/PXfbQHIaJozh74alOo5Z6zoyW/oAuX+omDUytiN7GM
lpPojE1JnfJEXbT76IC1anLzgXK2sqUH10vuLj0fd9I828MapKjh0xTR5AN1wxf7DsEEpwAPa7wb
7zxU5AyqYZsrFEymnhP+m3ccg+Mi7OcPjY5nY5flxRzOwMzH/s5P5QQd/Yxo38w6SOOHk9XzXSw8
5ZV5+8BtSYJfhNhq1MSB6x1rkLcNVBeh/nfc36a8UP3G8NF9MXQsenxEEPtQShtchtfCAXIMrAM9
OUDADpmDjrME0zfNV4Y8prrddB7Ilpxrgv4BojC87pl89V9EdhqbdhRCKp62L4hOJNoWPBFsP8rq
SZkxyJI4Pi34tGUUj1osgWd6Zb0Cp85DY+WtsVMYUEm+2il7N4CT47k6+EoSrlMW9dca+8Gfh9Jw
RysLDkA6rJvTNTUpfhV/Tgm8rz3GN6X6wFBjNacOVIjBo3S8PayWbIHG+ePdKxmJlA9KL/XUDsYv
Z/qlUAPBvzvhBOf/Dd5JU4Uf0Tf1XQaQ1bT22XkGStbiQuLuaeLcZVndiNYZ6xZjJhIz4CSqxIfF
S4vajvaTNnpqnfk7lgzqHZn0cCSq20uypxp1PmvPp6d2mvm1isqqlBCQX6x4gsFW2LtiWFVV5Hbz
aSpLcjXkBchwZjgX7xGX09WOJ1gtnznVmMZYQVTcLiLO/z6AObmsLvpfD7v7mFp/1+Pjv/T0df9/
8AndxO7bCoC/JlBYWvVS/8vlhCRwaforGmtkT5BFm1oeZDjp4alFJFGGds+NFpcsa8gEzDXTN/NU
sffOHlo0aHSkB4unumCL/5urNf//mKYvOucA3DdZKWXlZcvhAQrktNU0RWjTY/S9YDw4Uhj3TKrw
NLvuI9AO9bcszT4aDsdLkGfEpPSZDxhji05PLPVzkYkt6dCJhzy3NZH6UVYjuUmDbtjZhv/K0Lb0
UXK0QrES1ZZFRlmKFf+GjPlLlsnnlgkSL4074lkl+FQL2KJIASldzsLUlBx/hz794sCvbtYnMvO7
jtkUSB/bh1MZNvKUZtCd/li7XrID29p3c/I7i6oZzz2lxR6ZqUXA5N8mmpTLWZZjwE3vOFp6rKv/
oMnO6yjQzytwBtop7CXxA3cdWHzC+pIQO283568/5RO6SzznLnwNOga8B7h4DZd6F54fSsHiUP8h
uOZB6ySiPr8nEiFPcyduDYk5rt6l72tlTspACvyrj7MquIStIQ0POJnGNyp48Oubmen/aLGcbhq/
9hR8znD3YvqMTHIm8X+LvrLSfryL5a/KbEenk/1qov4VkYs/+DiGQzULrVm8DRg56huCW7ugNNYg
ZmD3axvQYfURyJ/9CpOqyqQay/SF5umuVQ/cDefyEnHD4Q3/3cSRJHKHNxCv9hCDYTLYe2W4TGuI
oslEfjprEWBp2fmgr8s9lchknBA49MkDsPwxXnLf7tUrQTWBN3OsFd1v1aheizRk9ZfY7AjIXK08
pYPhia1J9FGHd3O+pjyOT4GEjOqpnFLRlJw5Ekw78+oxaSvBkHBUrOt6FsjNEJO3cJfO8a7/s+mo
/grERWusWoXfQQBCBthwCYmQzMBFDPYyXl28h1PMaP93isdCwzO/lg3z2bfbYj2c+L87VtdPb/2i
U0pMb7Vm62mbq/wJym4i5Nk7bVeTV2B95A9ZuepvUnYasZ1t4N023bceRxEYS5WP/c+wu6oPGkmI
mTjuQXiO/pfEnCtb2PpU8HPslIkDx89wfSPyLcdkBnw0gVF4L2AIbyEX+8pwGM85boMFXWmn7N1z
MrdOCyEnfjLr2YkPcQn/6SKIEh7U0F5Dd8YuZ5I1z1ZwpvoRM//Nzw7WGhCLBrafhlkiXDOw0/Md
5jUFTynMM3+7MmwbtX6jqBVytrHHryo+hfB97wFllwdMp0XKA1I4+DizQoQP52g+Aqg6SRDwQAOj
VzAWN80GXgBtXmd7dt1cOZXav8RjeAIXO8rg4ZfcPEIrh20HljrVbTSeKMKQsp1h3KJSIiNojNNM
r8WtgcFiosNsufXkaYRmcpTk/tJdGvW4/1WTsuARHkqaj5TiRaSHbU99zN4LXeMIwrmr8u3Ijpmb
terkurdSrhxpR9V9mvvAynP2jHX/uU8gzUm/01zZYfk5gJTCVCkX/I+yWnHzXvTNVn24avrdLPrK
HC1a7ayoLHgWasuM0xEgl7nS/ItCOmut81qqeyxz6Jtc2PfI8PSZSPpBhJ7JCIChx6Wgz0UjReVk
Fwz0LpIwfsosyMgliNPi6ZqxsmPih9bTHa+FvCLkpqS1snDc2pS0Sa0wX1d9NnCePm9y5fl9VVUI
yNQ8lcKf6q78W7q+tugLuagWr5ypd4hfVT+pGTDo3uz6Md9q6dl8/lfwSROvHMPzR2iwB9/ZE57S
zyY4ua9M8f+kQ7gRnbV1MeNdSmQcgkG6CSSc37Ubf6Q2d2MUBmQlEGCQE44EK+QsqJfAu9byaYWp
Xj4wfVrtUSpWcmtqMBl9dv7KUFrHEm6YLalTd+tX7ujw63Iltq0CZZeGKx9S+SBBe/o3mUBOm1+u
WRFq/yv+ulKLp2/kyFceDpACB9L4+e6aGSa2y3sUuCW/m2LHFC4B0FXwERJEInrhRHmxsNKd4V04
2gY9WTo6fUyqVpV+BqA0/iAMsYt30IbHO7SbhEFm8UCXewq7Nwzj6ZnUthrSasAfAGMxL96WMrey
+9x3UfsmWTFeKdd2EvA1n0Eqdb9aZq8fMAdCF4nqMHgpFYCLJVGzesfLogrBEqEXyPSv/0NcsBWn
l6bMgPHxvg6nxa69b30pKO/mJHiOcL8bd/Sbz9VI/B6beH3ahI0rHCaZbjnv+W7T8m1mKhREI0I1
YjGRnQVMIokbFdYhLcVLoYU2dwX3pveXIARCg2Fn6d7FO/BZUix3FzFEuo9LwnlqCWiZOQqV8d2B
rLK5Mxvf1utv9ppSwTgQP5JziLsVpLTrFHtWlQByNO3TwW7PIC3ZQDJBmnVgBQu/dYhz53cZcPrw
GZ2hS3+a2Ov4T9/mTT32Ymqv7OGW8cQA2vBSCsUqX9qDDz3+1TFeeD9AuXXezTtH9DRg9u9qg/Dc
F0x4lkY0CXpsJPA5qs+X1JoKALeXs3FqhuV1o8To74ws8RPO9cTEGrvuAbO45Lbb+h1KpiZKkNZf
Llo+D1kcRI7RAhV0u+VSJhI34eYe0GJI+nRLq1qY1a3tJgYB5Lki+4lzjEw5k09e2p8ERV0EPJNB
MJqw91IAQPdFYPpqS1mq1gQT5kHt24hR/aF/k5A9z+hYSeuaP+MWPYn4UshmzzGCCEhTXSnd+plL
3ZTHzpjVefJN8+cjMPz4YGQqxw0eLTDHjuGtvo9IRCk5yGYlBIa2+lCdZrB1kZGS0u2iWpc75DZA
Y03d9eIHzirGR+ddxV14nnBPDZTUdJbII76hrL8I+cVsLZScce0RaeSFWv4aMQR2gxX/ToY7Gv90
m9l2YLt6yE4MP/4UuFqrCtul9yzCqWUXXopt28kcObMVOmNR6JuFXCNDsqtpyl0FYKgqQ4h46wnj
uppXb7McAQpLTo01NpZXRVrnEKPu3c+F/vMfFYJtiPMY7gUZcGPwC+A+1GJV0PYeIGCWN5Vdhx/8
pNdc/o+1m25OKWXx0tCMJuIHHql0iJQowIpj70wG6M+o/lgfGMhmC/w536i0k2U6l7BQrXCxozWN
77ad3fLrUgjgpSJum2MtkInVt0KY3dnxgiobRtVreX6OivOAmF+yAj/1h1j3V92tpsFtrxUwmF2Z
6JqzGu8Z/151v8dmrWdqF2g9Tz3DkCkTRnkacvQtK4Oq4/bANfWJc3MzxCyXOTXSqHln0PPl/itz
8Ed9Pzo61MjCbQvJciO6T0AU2tNXdEpJu7FiI1n28pnHGYX9risEBoME5kQEaVBk7+EoDZWta7+F
fAZYbCaqsdpPOqvHDigSkrq5vcemQXhlK+EhRzOMa2TGaKcyHnzHjlxyBtFG17pOJYov7wJufLEK
pMDTL4Fop/6JFFbSCYWWj1XheUbvGYoejOGIMiM3PoJlbaJ985+Qf/eVi/aaadgyTAlRBguXj4oU
0MWh/4YcNly2YG5PGQqJ/nQj55Myeb2yrr/tKQI+8Q6kVy9NMOQUvU8853iAwzaKuNpujmSVFzKB
q5Vtf8oH6oooLkYKPB0GFGDSYjyTMUkeiL4Rhiyjv4gMfiWCOhvvdew26CgIV2MobgZOGoSLc1ke
7kEObrwZBdXyvM/+R2JS1uENOpMb1xibuyBfFNxh2OCD+ok4ulGmiYIGuquu0vDkEKByB1DwDEOu
vbQumXsi+7P8RJmEMLJpMacLHkEGe+n8FIFq2fPEC8776sN+m8cY0HabDxk1ODmQJOA7aTCr43wP
e3Ld+6bd9uhtSU/MJUftLiWF0/1UHlWuZPatMtRJMfLRDNyTtwR47wA+XybS+f0F787FEYyqnaBn
MCgJAckwcJVk4svPNemgq4Yis7QkprSB4K83fMjxchispJzopa3hNPJbAdA2I3enl2mH8mEzTYSU
3HjUFqO4Iursw28PSpFDDSkwFFYsB/n8nhvmCttWOaYj1MPAg/4ldB3G7gJF0absbPkCSg2ocTmG
KgjIUvRjloBoiO7BRA17KuNUdP0KB3aoTwqmGrNNt6PTIDbLExfF2Kiy+J1E5nSYAukhr1sGjhUu
yDm8STev5yEtraw1ZL+T38V8XQ9eK59BOc+mrZObx+X3p+lydWeG8qFfXD+66MTVOLCDWORSxqVM
FrbHGmuH2QJCIaoqpNq31YtVA7x4GVyu3ov5aodRguaCZQObpDevBSJFVVlaTv7kwqu/Eryf+tnk
2eXlRjAyn0524N+W+C4kuaSZvROG8Exv61MhPgJegE3OSNBHXRPKYVfSGBlgNDr0p8B9NwaBm0+f
rHBR4NKJJmVOvBJNxI3Ga2JkByAItbQ5rJ7XxIP2xgbmJ5IUyGrpt487b4eaqFlGRthS0VgqV2QX
qOBvCoJgnCwgd1cpz6erWHrC3giESg4GVAcKwGdqi4Jgobll3AtZWBhtgUipQP378EKZSk8Z+gU7
QVaGDu8e+vGfDE3Kb5LnpLGcGefHrTdSfL8Sr43Frl/wZqJtj77Gf+rFp1RxltbjhwtBqI5q8YC1
ABBMukHtcoCPW4l/uWlgkARChagBnuzb/6cKHEelmZCydjpbg7YL4QksXSs8b9DzQ0boV3Kp0l45
GaHjaCL4m91XqI0+3VfFdoESWapO8LNDWkkpDcUWxZdEhfXPFNAnNk773GkJyz++2TMBLZBIdYvN
HQc4zfw8AdzF7mNXKj/ImMCBycEKex4RMwYAsMemyO/9glS5C2ABWyGKoD2BVAORM082lhn/MZSg
oiaOZXq6qK5lN/127acMuyXLJQ932bueGKz+R2/E7Fv3EHxsy1SyC2RibBykKP88ldggbdWDmWIJ
PJiQpBkVWEg0aHZV/d4VUduzLA67soHqmf6U+EwwEZuqfBlEQKwcEx5ZRXWTKrRAKUKmD2Fmij6P
GFv6mh3sUxanzYOOoEMtCNH4KXnbtYytZKDbVfRAHJ1w/FV9Xta5cJI7mS6k3XF8I18jrpIy0hE9
xzgnvz4PORgC2XhVUfG/YUhyNaNagFscM2tfuppLpDy4ebNILvuUv8UZMMfzyxLp6/+Ikg5vixM5
BU6IJ1ZPRdNfqbOFRDuVpzqzIfG0yir7TJFbtYeaXIEJsZdH3ArUyVIzDtH+ymumAteGL/J+pj6l
datuwkmjvuOiVtNazkZ8q1q7VNYwa8szb5RUTUc9UTwrjZXacNUVMEx30AQwmOX3W3IfgoZ2csnX
hAzMjKa8bxg2lNVxhJCDt6R60igC2Oi9+7jmmq3IwDFL6R/auqKtY/A+Wf81ifUi6M7N3ssHyMfA
teTJDvc8d0qUdz+xTEhg0ZWSFDdBRtTslp2lrzeJo1CXiyhuGesl1SG1fWYtaCknnBA0F7UMd98X
hMCXxA1M+sKhEKYfsgPkDlVbU6PTdowO5fAoO3JQRgq00n1cRpyEA+q5MF1LsT2mUN7ieUhrkGdK
eNEb+wYLiDV6hijwtw3bbNxFqSm87hvJYiqjwdkGrRFAXrjgF8WObYfNc4ceixZ7k+smSVQRRey4
uGxzw0CcbatMnZoq3c6PBu1DL5JuZN9+3Y24pQUleX9QQpgAZRH5Iq4H/8gFxyNUw3CbMOlxrqYO
dsoYFzTEZl0c6aqYZUiasLnpsmyhZUpprkO7cY8a8xlhSwvwRb/gmi1aOU8KuItaZnCFeagjghZb
Ii0P6RIRL0TDgtpLaxIVzOCmP0qlcVXGhTdtGve1fJcIiSC23bgoaPiETyWNS93NRdc8jyuhEOGg
lHgHqLsXD7Uu2SBmFtF0WZFXNjKU9WO8EdWw2lVyRaQb9NB2UhdLkzdPmfcBvJBwUU9DvkE/wHZJ
mty+HJULsqJKhWLddC+TtmZQnvZnoG7MS+QdEkkvbXDMkrkPEnTS4xzecP1uGU6I7cUaImFX7frf
YaURHP9lkVfriIOka7SxT3VetSdH4a0UO/WoO0fGUwcwqpKzKxuKMfpV73qLqNRD4kwaWkOkZC2P
oXqaoK3yv3+WwhJpn8NeVG1aAUaQ5W6OskwDNHMMcQIpji8y4Sb3tfU3XoKx25w5drOgvAzoBTfq
lTW9fdAvX9jhYlZvvEFBll/AooagQdVZwGsgk1JclRUCjCat/18LwDR3Bg5vZaFXKggSaPitgdG2
RsH3T5VSF+7C9BXJ3Lvn6xZ9Bw6+sgFFc70Qq6qlIo5oGiHzYxrufN1joFJ5VTHKHjjpp9WeQy4/
64owhY0c5hA8hasFje79Qm950NFYcwf6aO1lJwDXymFl/+bkJNEdhAHh5+9WGIqMU9oXjXHN6n+w
9faCB8gsOudzpq8d0yTMKMR5rtaBAgIoPRqC3GFBUuvdyNgT4IuxrZVQhh5ramWAeLWQCZWA+JKs
FddBXTLgw8oVXos6nlfyamAheAjSYRHouR70jcqyxqpKNYxiNdM1IbYxxGRB+UObC1jlzAA7O5Lm
gJ3mGBYG2d4X0z2GERUiO42EUrVL9e+gUnBPWsAO4QZ7xn7li1FOQe5X6RJ1Cz5rggg6LGtSrvHt
IbGGdC9vIsWeZUSKL0ejy934JoOzEZ9NjcidNX7EBe1KdZLpdbsxIkJjgkb70hskJjOZYMQ87H7A
JvYyuqkU8k9/PTt+t9R8Y2CYYNvVSUyMJsFVML7jBXAq4J0D9oMtA90N+aw8w3CGfkzoN/+Gsn5U
1X58z5bvFc2cyW8111CYEU0eXZ20OLA4rc6TjZs3cT/UJ3HSY6SiKWPiaIOxgSbfvttoZ2PKWXUm
bjgVB//+a0E7Uv+XjICfO7aS/n6Zyb2rENzlmz8qV0s7sRG5ypWHf5nQCvPL8pB742kTqrU4elvd
WgkQWMfsFq8Ik3CsJgJzNR/p09MGqSa+vyRiQ6NzDfPitTNQq+Iqixzi6IQJuUexJK+OQrmdXuZl
znGMz3vRMS+9M0s3eCBMAeC2RjASNB8Y9JqNOnW4wi5aPOpwamalREUKr0eIBC0yUH2z5EyYsVyy
VbRB/tbOvrqCHBlZc1msnw2m3po5mnbnD5IPeZj1zwnE2xqtEaiVk2RSq+G3Ci2iqvYoPyR2qZwy
tuMorsevBHjc8WrOLzvCYGCE7YmhnecDYPeeX7DdrWTzfrhNE8YxHDB3AEn8+Fx6MhUPeuFpxXMx
53ZIjUrx5AOgAWRxTQqkiRYYbqmpj3/YIHGKnj41/xxNdTOST4+ZeA1wh74wCJggkf5xbQw7iJRd
BEQQ21dn9/LQzFEPUjv2f1bGSzXEgKKJMITZHBe+KHR9uUXxiBZ6RigxAtl80+0vu4c454nyrtcr
IOCE5njZXzluBEi8F86ExMA4XTKf+euUQB+N8XFIx5XsWjnPVrcG3OtQOfyIe/Ts/V8/VJoyj60a
HmVSEkWN6Jp4NSnbupV3x6KKtRo+wRqE6DaG0ySFHS6hjCWmCwbcY1tyDbkZplyZurS5s4xzjyj4
8hlYLxjusLseZWHq8OWMvYB3jXTlghY1SswuuReFovsgBR+SK/aGo7jtit7rRcx1yeOaFUPdAvCG
gumc8OtUsCkoJ2dt1Ns8e6KRxXl0RZAE28sIaHsJ5yxJJxDOvyYJDk2SalJFdxcqJFXSvqGbTBJc
fS7yMvPyzoJVRmtVr7r4RxA7+5o8uNTZT4OtLHLXU9FqTXvKNODa/BpPsx+fnfwiQj/5KP/V0EFK
2vWYa4k2XGmroBLznnDFNk+lxGLB0JaFvLO7Rgs6IH17X9VRc3KBGkCJdYgFFEsF9uldHPNECr8n
Of1U1KRINt5xZUGlSaLsYMy+XWueNSrwrb6hZjc2kUV607b8DjRQVbMCUDaiPkdf8IaU5YFaZrPn
E1EAx8+la1YjvNd9qP0J0q79YDvOUcXVjLtXPvqSllixRx4gR/RCIT5bw12yBl9PbCX+T8Gp2NUq
mnYCt85UEcaodSxP97D9PviJu6nDbI7F6DkD6L2GgtUMzgf6qLxMTavLg3PshAmWU+ZotKJeUfFX
cLpjZf5Z0Twl2eNXaDei2Od+XPGPUMuj6e7oyjVyYQV6I2uHyuhU8IQZOirNXBElHlEqfQ2ZYO9Z
QIyB3pdyPx0jo8kWK3Bv0Fd1qUK7FAp0XIMmOHhrBmKtUwMlPshzIyRNYDuZyy7Iu+mwgf525nN1
zdyomBhiCYhccm81JoXhYgBVVk0pT9xXUf03E/7Di6Y1XPAG6hL+oAePtt2kmyb94+JgRdYDdibA
+5/iWTnPkaQ9Mw/4FqxoXDeiTW8kr39QPBs5VOfzuSwVdj6d7U6bie2f+wQSAOWp8mFCr2ZFN/Yp
aPsrs365Qr4fFWtmJmaLjBxRm8c8TWx5tTpUwgdvO0l2AJMbr9F3ubyv+ZlBrmoixLRctSWM7NYf
UbHcpBsvzW9UYUeFgg2qklg/6lixaK1C1TBdB0FN2a9HZKsEo5uUKFGHig2aL8wCnB94EuZbMDuj
oL2aQmppCrviJKgoMeAWWpSuKsbkntzvjo3udg5wfAlFomoyFqtsn4/cEiPIQJnMf6vgpPTO3IuB
o3Up5HaZfxwkG1ZdmuvyItcBozUn23/YhSjSIW7wETex8ZX4fctLWQ7rBoF9+oOoWjl8d6qGCygW
GI7kvsLYAuSYy/QTMnadtsu2DVh4Yg4QSeRckAcxn4jKFd+islRrdEyeZafj3b0Gug2gOw3iPCRd
hGMS54o4FW8dPk6vYcagSZc5MFVLsyoY2O7aLRiZWaLJdZIQ42mObQrh48qVXzIMqTRG0ak7ZUpw
Kdop0v5E+T4V2UGr7NQQ5gTB00N0RjiONrrnQ31Aa9CRkJmgoa5R9rqA46mdtHIs5R5sY4qpKuSA
gUJylMkz6mp5o3CCxW2bXotLrC6hW4x6AtVyt1sdaqXN6/OT5d4PrVAt7u3JISHFfhcHF0DoYQ/a
HzV59a3vyNycMWfNL0eI5ifqSL81u+yZ8GNCVIwxtWW426zhETa7O056WEX9xn7Bov2DEjkolaE1
rmgQFN3HIe2PVbXXvYhyJQogbyQon8HpMwxCwplpTI3RD2WIPxPz+8W0TYSqjtdZWSX2Ro+y+KQZ
2Bs5AbrKwDuVWHEmOqh2RRqJK8o9B01etHib7Ujgo6TRfpK2WTpQjRJpM45+OHNcNhtQltBcqq9a
l6/IIr8u0drrJep4kA/iWwOsw+eVFeZtP8e5YywZeiwAvWl44upBn8+EK6aB9qNE7Y6km+TkJl+X
N66xPWJweyyW8iXzlU2I3Ln+BXgg7m2lA4szzxQghtAXRbB8Y0KnmHjWZDmwZIiMd9wERFzs0q63
StUBIID5FZUTqrP4lcNhRSKrRvsPwr8GAGkF0bMB3f6LKM15zi/dYXikTGhKb/tcQbozDJG+VHu3
GqLFVHiuQCTOe0Wss/nvge4o7n8BO7xSg1pgvw34JsSqVTnSIb+i+Q3MOdHycllW96gXWLIT0XCm
AKdUTrJZE/E8EFjm1i17G4dKEuVKXBJkdekRfSFhmRCBvicH8MF6mhYoGIPMnft7lHXdjtGJC2CZ
QqJmk6B24CEVzsz4koHzqkTg4gvVsGjby+BRoDnxNDU2Vu2vqc7a/wf7w8vWqCvF6uOBi6ynmDp2
ZHDiIujHsiFTrLUQStSLYf72JeNFmLSD65HCZnE9tixPUkuDTC/CVkA0xPwo25i66gOQwNw2mU9I
Nl7v0dnjpR/QXEw8KNOZ0KJutwhsMD3/7IFPRJjewGpGxacJcSoxVjU8c69xlliYY9jpumUnVEci
IjvaGYjhXsPRyLDsiCJbo9MKr9PqmjyE31baNdZQvfCMq/hggKjD/Vtu2LGLSBB6iFmonuyaZ/ll
NIfHQPSeXFWS1N7IdH88TbOieJCuNS9dPTx5vCZUosbyOF4OMRzHYX7T1albWARriSg2i2MnvwM6
jMqmsxZbOBJ83RMITlUWr/1aeohSqL51oIDMKKSyOwr2LTDbCJVJu35EmkEBmdqiJMrh3ecYHpSr
EuS0u7ZMvOOQr4Z/R6DEEuBfqYgq3RyRDI09iRA6W5UZczNl0z7SvaOw1itrHVSxZESAuwzjRXxn
L9QkHYpsXuTVM0LtSdM22AzS9t7jEhGxmKUmO65Cb2XwBZwfxS02eX18gucBu4gHAzHxGF2CxLzE
1srIJnoaCIFI8h5GzWKLmgQMDLu42qsu4qejvEmsHCe0xSvDBpEq9Q/MaUUUo7EdJY7d4g+gUuNL
GHqQaUCt1B6CqCCGXs/+vagc49XsLl2dx61TlLEDg4VaIAyCrZJ7AiALjziNelP51G2R2jWku0it
BEfCpiHiwQnxbZLnKSYpRSW4cW9QkBqX+l2qyuuN7sxUZRkma0nIsok69kl6+OYRRRbxeVq/BMU/
c8ui+TFj5J8Gle3nAYAyuNwyGpn//8HcRdxw4S9tJUcrbQFJa3adqiN35O+YYliYfRfpGx8mHhTP
iumdrJBEawDqp2yagPhWWv7gvQ10KwhlddGHwBnLtGQvHBVDH3pH/sZB9y8tBTu/GkNgefAlazV3
lz81SKFQBBgfiVFXZ0r0TBDn5Q5lm3VrY3EhEb1sJZpMxxaHcPvil8wh2V6fumurrOeU7QwTpOMl
cs01nhYOFoXf2bPNw8pgbyRK3aw2viDZFBpDldw0m3gagfjeerijXEpA2FgMTaJskEavipr30P7Y
no/Fjzbe45fzJVtmesIw8TWvaaXQ3c0w3HnQnWzipzNyQh2WWTdgWleD4o5JpDfQ6Wd0ZC0Oyg9i
/CMR2o3fb7exahIBtxcTlf0LWoJpYDfQpFNLtHNaNPioW10fnxBFXHBN0kcqe8/U8GlqmSs8NPGD
J60SwIWbDqHsZ7kLpUaCv5/mAev1FyEypyCDuuf/PYwAJYIvJHfiDneMWpuVFolOtqgErxaD3UGi
JJrj63TWE8pRY9zkeS/sWhlGRZxKNQTNJYSC0WetF8x985tAJuc+iqQqoFSMixgUh67hJfSX65gg
uNzhMW/8vkak8pOZxe5R8IWRua3jF+qI3IIeLeBp7+OvV1XY0v+DtYzOHGv/CU0FXFrqEhGAOGr1
OtGfiY2IXf95UZwkiDLTVi05jVMDHsh0luP4KeQ5TDKg/3s+j4ujOUxMJXFGG1VGuHdY37R3NLXO
rwJD/mjrMwJxSwZMeP0lw2ZcGKaCWkVKGlMEXvvtckJbQ/R6hmFcO3SEuXaJCz0UPyY3xFQcm4/2
CtV/LiENid+PrW/Rt8YN2nue53/ptACv75yxdrWMwMIEeSxGciaPDr1bGvXt5yKpWa58eP7CSdpX
8d3PgXoNc8TPg8cpspepcUFOfwzbNsRaLc1kS55EzC6YBuMARFkCuBy7lQlyKdPY3eGcG1NXIaaR
Wl9JLXodnKcDLcHP6oq/zU/FEgSLQI9rXAUcEpLvikt6jN0aGzTYc5iVGwkmjSh5LFIc3dPsuFT1
NngYu4zHunD4Z1nxCcypWcjg3tonI9X8u12TgdCJR6sTDf9M1KxivF8xOrARIPjJNtxUBaSkH5TU
XptQQSJ53UULr3y0HbXrltA2fnA3S4gn3E6p9LAww/kL7BPeZxvvSMSDO1NKWbI5CkvQ+MsqKHhp
pv5qh0x8lAJb95GZJjwVwZZ11XBjtu45okYkS5dxUDXI+EAqmg4gOPQKZQjzHzQC3x2Du5M/mnUh
K/SgNtiOQGy+xFTbYdJ1uKbvbnLXk+c7ag5pIe16uYyebng5reeBr01z5bhSTvmDPRmUZ7banNHG
Rq/lZ/oD988kIzDQyfXTHKCtfgdau0ILSOEic74/SjQzf6dw7jz32/4T7Jo1nzErUrnGlncP1M54
XaVGP/sIuorl2j/l6a3EGVkg1Qo9GkZqSXJ//eIM1CNyuxiU3vu8hA4oxfILwOXYsas3oVE7DvwU
oA5bpFZWrAN/eU4nxBbovwsiFpPU5CyLZYh0N7m7kkFeRvwuUuImfYx5TFeAPCaR3248DlCeTNhS
wUHvNbNUKham6u9xkASUl4gNWJC8eCN3DN2e93VLis4pfFLeJiAqa33XlQCaO5ByxzN3psDgUoIG
VpeIB+NukeiIfWB8L5KtI7uRB/AP6JAcFFk3ZHJ7JhNl61VLVwRNjBpWWFX2tKYP3sUh3hvqzipD
pTQZturWg1AHjqAkbas/FiGEtSO0BMa+3tTfpDKSnoifdXQ2wqzbp8zftJ6+ql311qn9WV5TN/wa
+3zWSaAhJ4XgM4cZSo+iLmpba33uy2gAEaBvotGXGqprrmXQbk28/Nt+CVbzaUMsftmsnkisvCIY
AVlp9cn+6HUN9QpkUGRByjX2velZPfzheUYNL1exholXVRhqXLgGvLWD6Wmn9PkuypdIlYgn4iFp
4aD73EeVgGs/fBynek0JIomk9GZZ9AJDFGoBmEJ2UZ+sKp+DrlGpb3yXPllqAHTf6JuE/tx6JYEh
3bKt8ztXiHU68Qi54lRJZ+VSSMTzINUCAkNYL6tw7VG7LIEb//BmS4L9IXsDLvRSLG/D5xuDJaxe
F2G0VtywA18q1bKQn5+eaiNNFxvvyQtJY1WTjnHG7J5IeHzrNH9BG1qA64xGoxBeSK/sgw9B4TCE
05dB1Ph8li5CNVoT8ITOK0YhEmsRBNMBM5nLO7v8QKSbQtON/V6dKrDwfu4Iv18fu3j/ynuzPTni
TYz3hcgP40nMxNC2MytQkIYig8fxwmSmJmJNL015JbRogxkmPokhInRx0LAHhuTxckGN9aLLepqr
kq4MmWI4QYxq/0VX/0fuE5ExEoKa+BZMiyDXA1UBNVZUYUhtX1KYPA7g39qkvfwer/pmfNaBPXT7
eOmoT9T5I1nW2sms6eq4PXc8kwOBmcrtDcPraFfLJ24pXuNUtcFUPJX7MyIgxfEtZ86LkSgOh3B8
anLIhfpZIe9akDQNlImv1VxXdTLuwfnUdARgU8+TrGG3EZeXRHrhD2zkgEFiX4TORo8c0nrmk9Er
VrKm2oH4TLN5ytUBvymrQW9lfcmSrt2Y754HASAXyi0VrvFtXUHFZbG9x5WR/k6vyCKkQPMxNCpn
r4uujIn0RkkzzBR9PWNnkSdaELE1V34Shl8I4IITRSOTzDSi6c2IbulwhVNOnTz2NpLGjTx27uM1
f2FCTMmEEynvGdYj3T6ahB1ln4SySrAgO8GT2q6+Cwas6VNx8mnKC9WNvdyXotbAi8QtdBXZwxGU
Yrkk8lsLrH5Vs0dFPJGMQw98qpxPdcuoYDV5VHksrqYlzpTAb9qeagKIKnig8aZxz1xolinIWhuV
OSQckCU7yDNr6mfKZWAIfw+I4IG9cuy7uIJrlMV4CyjZk0l5rn4qtODeMe9fzkvhUiGNRQmD0q+2
LfhU1QwVwkGssmQHBdBvDrxp7frjJzdzRWGG+UIFRSTwJ38zAKXWD7SJVj9hN15CEuj+7savbpda
JYN2zJ+R4CMeJx030S20PcmxU54o8fdYqNpvxOPD3nesiHLWETzp/5VEiRSycqmduzaCdDb00CxF
d+0w/3vJWS9JN0u1L5KbGAate7WXU8auI0vaNDisaT6a2miYxBtkj2ldOEBtGRgOVzQRYMs32Wdf
Llz4QRtt5vvUcD7DMmAmrpdi4ww8VPKCJMPkUqc5nV9LQ4Kd7WNOkIEDCMl2c3RlnqUG97PuheFV
0Xj1G3TiUoVCdVF6oG0ug5y7AqG+nQpawQREnM+Ta8IjgKU8EDmYR0Fx9BtabM+tmi6vWe6r7PUp
NSpclYQtdk43vlENXnkFJgNubVvJff+t8jtyAqpUsPMg2uQcG4ta5lQq4FZyTaRXi9AQINbPf3XF
NeCi7zSxUSarJTAJmya0VAYaUIbbMVgN5Kdq3ql518+lnPAZs/HDLSBQCzERzDsS52kWr2O12SUc
p1jxZwBCgPRmFCUBfO5deJPw4XWy+lNuxjcAIyH6SoUOGtzTFRPVdq9aju2yov+X2WM3kBFAtOtO
2VWzkb+50yIUIZoWcP5ecE8k68+dNTRM6CpO39YuDdOTXM/DMcJ7G+SZo4oOve97W+Ug2LamZaPm
caJoxThpE5c64v/kT+NJ3+wpTy1FbIEX1zqBbVpE2GD1++YtVSLFV9S2q4kjFrYuDr+2krWL6jef
OYuGHNuvxby4rlLpmXqrafOhBIRIE2jNwjD/IjrxlHGBIw4iqE7FTQ++jUZ67f1UuU9Tc9aHqfky
GCtvPkbz0QmRWvuh5he2tPHXEgENAPhsBKoTb+Mvq6A7S4V31FXSN+V8CXu1x+/J0U4pVRS6X8oz
FiXcxUmjoO4gc4iiJBzT1sINifnyzMaqCgtGHmtlQQokGSBXK4zUB73B9Qy3aZJ4AjBf3rwJBkPf
H5kXwYMQU3ENy05SQQ1JQKWUb9nVdke5Il2/du5q/8shNy/h/qaUHunU6X+RibsX9aPNzQk8b7MK
cBfrr+x/tB08M3rOd903wIZe0Rybyjzhl2yPCPPbtmJSoB1wT0d+fpd4I36+Dnr3aco1vhUYPYnP
3KR7L33Iee671je7X+eV5tE0dPCn6LkfZtFFSvHlAuKg70w3xiKnr2N/+1pCfsZQ2/VHYzjibOpH
gl0E6g84rAUqFaDY0CcOGGcrtYa6JZJeTHAN4WyBByYFO20JGfr4UPRNPScKk8SNNGbPKoxB8EBL
y3P8EmFjbqcc8+xvZjsif3J94nFyx8ufjHrZFc3Js90K+wWuHW0ewfQw1NWm0nJAkb2njUvZbhc1
fbX27q1YvMgKulI2/q+e5cDiguXysAHjGOp2RAlSyJSS9NuVCTHPv9li6CWE2rDNcZAPzZbB0YdA
I3kz99SvQQyo8YMCPsdcZjJhsX/g06x8RYO3onqxAz+7tB5QXB+D/UeZFraw1c1nTONAZQA6+aax
6eEsfLP/YEPhk8PeVX6rU0p8Hl/Fu8LQGIyeHB6oINNjCMfCCZT4hsDJifX1gLUwn4duFnfKsHsy
026lBllMKU5PiSAzOVHu6VfsX+Swnl5RbTQGXydM8aUA3Qb84RfoAcSu/xEobqWP4MiWg6fxMbYg
gPkkFlOobiOACyQ2VmGaFnM5lUOy4V6LUwnir1FbZb1r/k3jEwCMUXcDqOCN0lvHOoCmAQP4ECBc
IDGJfkwL0o+oOY8874xiWUlBk67dDDxYiBkuXRz0SDaafXZQ5OSulONIIqCdcfLlE4QfpqTY3pR1
Pi4SnxVgInQE1cuwH08r8UzWPhTsDqXEPugDtmyE0VhKb9g8oGL4aXXStvUnY9/Kcv27IaFUNfs/
ZfJ0mKmZCK/zRtyW7iw6bM6kL4BZOy+YlqkFFlZuB/sa4q3bQbRyMy8qs06TowLwf2k0ILFi//ed
z4AsHXoLkswEQoLZATjswJ7HMshHeao6rvIMc9e92BTRYpySakyfoBVPnW02ZreSjpZwmZR6mo09
q6tJKEfjPft+Nt3gphH30H9ItVrV4o3rIhc2fQcVWTYc5ZEixC5cKDS2RiQ6D6iXRTgE8weKzV5a
iUVzk2rHQgRZc9t3yLsJ/7Bx4eBM7l0LCseq6voPb58Tq2Wr3QKreGEKue7MF99R/8VdkcZ2/mZW
Qj1Y1uQgJwDTE+atIqslRlgAsLVLY4XLspodT47fx/t+O6funAw9iTCY2pK3Ps657banCV8FhstJ
12rWqu6U4M7oBBe3sUsD4SELcYt0B1i3wycieJCjoiZ1/NUuHKFTOjmSfnK+Fs0VsECGZO1U1RE7
BxaDX+6UrMZyHtoj4xqT+EQmCazvMAEFGMWwdsWTgtbnBy0OMo7rHERecAECJ3nvYoIlNA/2t3Am
lYkrWTBvWXf5+4jbNQ3FMAxlybD/7q5RL0lvGTkvRz3JDP1u3xWVAL2CVeBLQol9B1Cg3jTu6CNs
XgemwLbqp0TbB3VNROP6y5pf85nCzR4hvVx8i91IPZ4unDja57LKPQ74QAOIDyNHCYfwQ7DlEwHx
VyTwjjVwi9a+bdFi88oS0JFgh+UsoxfCnHJeKkBN8/5qEu/WG3SMzPhFfZYUaV5mkFWU8iQy+wEI
tA4uE2ziYSprhv8W9fBYJu2TljL59fMiyTcJf2zaQ++WNEsp0PmipZSqJKkGPxVcY0O67pC2f/b+
/brirv5rFRCv3ArEutFAVHAPEUXi+DeMyGp2863NSWlGBrGweGr8egGMt3jTSLZ8nvcsLds48waI
U4zc4X9IR/zV/DTZlBIgMpdjT48wKjy8EGTbLW8oMcDksW2rbvKy+ygtLbs4w96vYjW+vi943gTQ
60wK6GHTH3p6yoNhR4sdiv9s23IxesxGB9WdaIC0Hlcb6j98QysFjfCeKERhLdYthwJDePxtjOOV
hHtO7ppNIHOivAqwOEUFg+B/8y+9w5SSyEQ5nuQtij8n/jqGFyHWq+NI9apbXV5/NGLycyJnkN/5
GrhiCgKpPIKcVu0/6PpIAqbY5u0SC5ThMafPNlcn1Sh7YozNdh/PS7U3fTo5U9eOiT3xJFo0ZUKo
v7+JU5ocd+sPH7ilx6YbXDsAaqSZPAZUuCZrKKgsIh5WYzNmtQADdmuz19UcCiciWcioGl2cUQDb
R8nuDJFsSMmRtuiH2ah49Oo3hP4yX6zrpgqbvkP41r4UKuKUnDsLTBznqSF2zd/33jBjJVSU7AO7
zVW9P1wCw+sgz7Jjd49qd/dG67Yd2D4svEd7OfmmreLtYvR2HT0QcyH0ZnFbLqPYs4U9TF/dn5IV
IotDBu7ufYsVbEwUl3BzKU5JM9ssyby3FX1U1N4PXH0UqZIwQJgz1RPUKjk80b3hPYTBJl+Wo1cC
2wNBBSPR5+gNx+M7Mf5bqU4dMJxSd7HSPbhAbjLa+V5zxmiEG+MhQL79zMMOJTk5X8+XOChwMl5Q
mECm/S+slHPmMwe5Jcu4ntMj0a+duAYygXOob613K3Eo81uW20dn2a1HL8AAuebEYQTlPJuIcvva
FJZ3IGj2Zkltxn9fcj2RAzToFAzyuUEzBNK03gj7nx7SES3eDZlGpoIZ4yXJgR2qHdsWLp7Ys7Zy
6Ij9EZcD172juvK3h4Gp7ql+ap/JYLKc3OoXzJJ68TCuarQLzrOFFMYs8EPiNc2jc3kS86Hlji+E
l4SOcbu/mMv5r3Ck3e2KK7C/IXMV4kzAYwua7/W7EIY+/hagO8GJFXDFzGOHxRS4T6nXJzVKAmj9
6vakPUDol9maFtJGrb9CIsn52N6UZv8ujCmGu8rSyrzLlP1l1sz3yHuIvrpeSFOCFIGRbU9kELxw
HXmNT3IAIAD7DbVMXgn6m37jJlKRJbdBrZ6H9RN7vQMZ5/doO/f84+jjc108SIeC5k4fV55U4jML
jUD+90v7/1PHtyF2fayb+ZktjZblkU3RjZWuoRNyPr0fZxeBxgp5khBQ44vyZsBDGwH0ifXuqFP4
KfVpysStZ9/D6/5HLIdfcO6gCCvof752bMqJ6N92S5nvYJGPlFVRDBLg/3byuZVlWxnfTFfXfqk8
BzUY98vXgekjga0Jok99QWoRp81Utdbxx59x1J08hH9I8fMlxeP/7vSJczeECdljEsB8YiEYZM7S
fNFrQzaRUY4XmBRGS/zJNtX4k/xwE2Bn/OijvWTxNiRZ/kr6f4V1ZlWEn1YAdCfKf+b/RYi81m32
iic7Y3ZUIhgg0rzzpLKmRDFUKOVYmrrggLaS7u9RwENZpjc71EQC0tzJZveCRuWCwraAnvSGRual
fvaRJsez4pvr/IpU1p3NOwbzbwL7e5ochnIn1KAji7dxOkVTXuhqBU/EVQPQK+MoRxvKzN/t+K/q
ea/ELQ8GAynIqm+0N9BNgnaRGH0UclrfIpzPshY8YmZRZj2OLN1I3LT8CDqr/ny7GKAHo95Z2Hhi
AKV42URd2LRT6/i2X+O70wKdxxijPD4s3GyO0lJEEEXm48VNc0FNwcOZipUa5jQqLmSpHSte/L6l
ERyQcK8XPSSwsyQiT2o8xUsiamT+pbK5KDbmM+kdUg3y1K5whlov4R4T6OkZvIK0GsqDz3uB2rmM
A8aGOCr32lj8YoH+3fMBWt/cBJcomnvpxiwhlq/05THkQ/qfS/Hit4Er2FWOoNdiyZgEe/VkGeJo
fWZ821lpi3n1FB3rGbLxF1KMPJJODC3FZ7iuZqxQm/PIrKPb07//pljO4c63dbWZcWStg9JBElx7
gvhIn37msgvGXL02JX1fAJtmQXzgV1l/rsawTygoH3UkSApzro6r3gmIIrV/wDT+nSLZbkrQH/LT
cze1RapLdsZTT6ReDbWIvDEBmQ9ddoiSQkqcXMQ4OFLuvLsyjUKWk4N4ztFKSm38tcYaVabrktBW
IuuBepLW87az3W+ow8cyVfw/wHScWAYYPL5vco0hCz4GR7lInTukiJo3bGEU9fo5qujdxxUuAbxq
M5Wbzh3K6yFSwWFfVmZL3EMt5mhkm5JDXww25LjxPuhg/NwbW9f5QhFefnPC6M77dlOYyVjTswUg
NOy0t7IB9gSOC/4GbU8m+vFad6SEMaiCTelaGot6bkf11Td+2FB4/h5NZN+WrNdTbd7iGtyE68jO
2qDkLa8QuGQRH+7P19KVP1iRV2tl4lBN4hFkxlu1dNaf++AAjjCcWT3fDdb3EofJ0pALkwy5huiW
04g6gv/wAwtVYuEhtlAYO0kEHEmFXllsOdctfCrJT5rl9GjQ3yDtEKotXXtxjCY/fVVGUxZoxHvq
pepyvsZ7TUocEFGZg9P7x2ssZuCEmIGXqUUVk5eKMn/dje6PbU1WYLLInwrVQ9gtGUefak64Tfe5
v85GTL/99//1m6yErahNRCDGS93d6om/OEGjfPJFkJOUr3AVrxLnBRZhJAkfR5H6Fhxx34h8178x
KSWaF4OyBbDKQBEi6qGB5kQrG1vayVSw17v2JTGodMwkLZ4WwZJhz/RrbU5qim4bmpVpxq+53uBm
i6BhDxeAlWqBicg0TEVSEqtB17cFzAhUq9cxD3fx+GBo1vujLEauZ5qM8o8XKeEjwaAd4zD7pl3y
PE3tdGGWUy/DEc2hQCRY0mJ2WY3I/Ljr5i7EvsylKQPInINhXKGr1rz2c9oSkEiK09072Q2pu5z8
/DzKqiji+yg+C0eBPVs/xFutxA6DsNsCWB92UcTb7Sn7Fo2iE4rWSHWfa/XBVbVqgXmLplbFU53C
FWcKc3IDlA5xbeQgtYd2dJ8QdCKs5DCyTkY69PlHWbr2CFweIuDh23dMYwCh+a0QA33Bt/rZZ6Ru
8qnGb/xb7CoOqe7VlF+EUI6YFh5TlwuKULpLLz/ejOYlqBn8/ulWHYOoPfYP1L1krw9H/F20G0WR
DebPepWeDuitpDlGqzrfZOfVroMJU3ekWbu/u5pJdE18HHreO3WuTB1/61NEt/25dUsttlRhJqKL
qmSs8ZC11p2dtmQeulzIGNIolcDoTroUwOwdWcAIdVhp2PvkYJricRQvKR8R8S9AEh3RDWYZTwQ+
8FaigHogdjEvWxFIqmIY5CXIaCHay30Z0Khjwl1ASBZlQfD7BV0mcTPQ7nkClORaW3L1zoapMC1t
WSvpI/nLjAMrh59SKSGZkP+vqSOFqZNWjb0z/v6LCvdy3d4PK0ItZdXaAz7cjKLSWszGWhEnL0NM
j/5ui2qFs0WZ78x/IDMKxtcHbKVkZgYKFBWzD1Y3ov4TNqGXW2MT4mVxbI7hwuE8rZqx3EgbXgk3
9VU7NK4bEuYIVgWWwLCPTVICNk5t4z418GM3hw9SH4LhUXfaN3nhNJyp6TJb03Q1FUGIZ2AXDOud
t/O7B0H/n7SKrioNXXjSNFBRcvYea9UJKzonRvanj/Tu1mF2pT7CyGAwlf4JT+qSVcOE6HJznu3G
ykGVTTUOVTpOkkPs9FpBWidil8AELkUmHQ+XzQXGsMEvjq1BsZOHjMfvfusYQnfiFc61w5visS6w
06FCtXawllRh3JBtrRBJWbn4cd1VlbdzyNFslbgSc8SL0f+ih//7ayCOLZIuFiM0P6tms67UqCTW
Xc6jhucp7qCiPR9OBxcNOM1wszNppuS3LnNQgkh2t4kXPF1L5oR7In/0uX+lwG7VFFgraxV+iwxl
1DUAypOUFh9FgkInJ73eW6AimyzHdYM46U60WKCVY02eBVCvnwofs9RycIyEoyoIksKgtsSk0sLz
mh5doIhpmqphag/5GhX9Gll3tPOH+SWCEymnSOUHS8AuylnWmfJ+EehXzQdjf9C3FxqGTC4q3LpW
1bb1ToskkW12sOBIWDvbT+U1EevUBJji0N/D2kydXBwedVEV/Ni1RGmneJapkRSa4jYE/RQy/Cau
Tgm28cGJcYoZLxO4nqXxl+vS4xxNsSrGKAqMgbXiv1wZHftTKmuJnbUTRZTFgs2b7TNXdofzsSre
CxY2O5TSVoyNT4aPRDDoY1PFbaDfTBDimwJ+r/hZuLN8tKtxLlw+kCj0+xiaCEYBUwc/HOfRPxgi
fREZQqOpIBv5A//4yk1iCQ5uyn2ErFaJoZWFDmE/xpwUESCRRwhiSo2rLRWLg6tr/Gvo5qYjchhH
9MZNOaeCdr/e1JLHkn3U8B3feb9UlPXtjI3722Rw5Q6sUMqnnE3IZcoAQn3gb9Z6rmD2r7PRINPG
nhUp+hKR/3NwazN050O9En1ohhBW1QZZMOkttNTxOhqyxRRuElm5Rnb34vWdCMj5vuInQapbvqSu
dJLZmNbV2sKkuI6MuC/zMp33I7AIoR675JjAOwPgUxJlyzqdKfVc14kFO+1kpmbr0BdiE8WgzYTx
j9e96ifbNqs8vILY/6sQR0EfJU3G6fHSOG8BQK2zdvsOvlIsFTl7BnYrybSWzOKbGEarInJzeDcy
Wld5KlpmzaPRkLieGgnlV0TeRu5+sLp2dCz+vaZYUvE7cu+nhDu/tWYLRcJR81u1LUoQO5/K8XE5
TwDxvCFbKR1I57f3iZMqbqnbZBX99lzkkxpVqc3Gf3pFt5E/Myfv8AtUfEp/sXdO6uBwht5JqZj2
dHjVJCbt9u14hhZRS925ubfHZ8rTjbS2lmCByGEVZCP48A/JSC2zhO8X0lr7PvaDRFFqA7kSDdfT
dKLRmN7bh9RPdcIyQ45SH+ddSKflsxmmCRAJly9RtqTO/HfK5uLhI6/O0pttI4SiEoJ+C/fL5oWx
ineuMaQYgn9Mc+0gx6Qn8FmbfwfZVTxIcwQF9c0G9Klo0B932LksHht21+CHeJ93tGSYlHiQ9NeQ
1GrsRCudnxeYMGd4+j486KE5ZvFwolNtDhUIM2hqmzn21H172BB+6S1Ndfh+ZitzMTXlIbszHg8r
/J+7Uii+tDtaGL4cc1cbbnPOixAHj3fjr5gkN7M+FLk8ffuNPj4kvgPquS7dx0PjXTkqAR8pMMlk
DyUZyCCVrfHU1wR2Kvka792dcQaYaNPb8vkwUSPfgKWR3Pez8CTGYNaOk3dcI9Z+/xECUVGc4xfN
J5vmyagUYt3PKye6kBmMLYzl7ffCMPI4SiuT2rh+qUkFwZrBoVfLg+86aLZOHSNq/1skCdfzVkly
uATpkCLM1fK/+KBxFVNb6mpUp9k9SuG5zN4VOs8+JGFF3UfrbiKh3iZ7QLS+KBTIZBAK10ND28sH
HZt8hALeZlxFG6GYBC/erj5WKcHKgsmFi8jWZhJFZfXOqq2CMFFZ6b2LgF70yZPyJ6qgcPZ3/Opl
JRo8TXmqt1vZVgo7ccuhWF0E0VheIVoy5achcpTDVQkBQeg/pZhZczwv0eVphW4pfm+WeoXQspRR
499VeXdQlqbtO1cprOiK1mNvAx93feuSVq6yqyv+DFpBD3fCS7+ZnsJ0F69wVh5tFORsBchVxI0X
s6ZkVsuhMmbQVNVlZ4gv9OGRSVlUvnNZ++F1+U4Fg3nyUdGlPd8069x409stDu2mDPmqH/tbjG96
KI5glHZZCQh5HVSxzCBIZUFCVg3wG8PS7xR4njW1r8HL94McED2KcUSecxUipDL2sVwxPTJX/W9S
RxVsu+8kMRFR/7Mib4ppVGvkPf3PaXNgbX+m6uZkX343qwJh0Hhw9dsp7McduC1mXSobTbkHhKRg
TL8V7cMPwzlWHA1XUeqi7DFTrGeHGOxYHLWsDiu8E9oNWxnb/2JAiCgL4nuh0jID7xPG6vefgdON
SzUv0z3XLBOtfiN47ejbCujgUsgE0V5mCBi0nJuudL3GFUXRI+u3wUVFVirqKCyghAhNCfAOIn6e
BzX4d2KPB76gDBU8t1QfSTha/hJbn4GeRUnISi9rWPYHNA9RyFRbprRM6IxzkgE9z40eTdTz4+wP
YjTDlyTLBVJDfWn+OrMqzv88R0ucIQBC2YIVfYqNNZ5ZVfSYA7kyEFeDxErwuPltg76mC8u8XJ1s
SjYfu8ee1QRWLTnUrV0cFbXt/ltQPX/pTyi956qVmU43ryscRVeNqOAwaFDrPrdBFVD14z0a949U
WWHUsBd9PnxTG4ZXwc1Sib+HMBXVoXfcQeInLwNQhrGPx5Z+bqYkFbfC+azCG4Nb/w8sLq4Fl40N
1w5fphiLMsleBGXMOzZrQBRuOKAXKnB2hEoPrFbrSNit+/ersyLqGZl8NyClYOkTLERDenKVE3np
+Tm2Rc0/o5y2Z8nEk+ika20U4VPOehsJ5z2xTWSqb3wpSA/JnGSdMRtJDioOWEPgwShQGm02hM0z
Jy4v5VyeAGnQruOgDop8KrQOaZ4hs2ANK6TOmPgw9tYnD7pGP5HbXwR3EWyUjLywUSpAK299Fcla
3ymhxvRI+27nO4MHK1/SwIiZEfUkZ3+5pn9ZIgKyNfoS7/VjzcikKTjzJ+C32u14XoPKuLvKecn1
SUyQN2zMczpTWZWastcssDPIdOSgrMXucOEj+7MX4ZKZc+EiONYIRP/eeH1RszaiJmn46ADlEuWC
PPjY6h+jaMTP3vmnOXm7kitz69Xv85xxPJthKy64/spNEdHz+2wudkbJkMNcJs5pqcSaYy84ka1Y
bdvZs3zrFIS7UvEBvELCi8AtObV/4hml3tXGpeoo3lHFbPG3OKefois0jk7EryQ8kOHiHbqWkrRR
fc5yo2VffeZSTzawHb/4OkFItTtmYcA1pSKEIJxTWtIXfQqiGqGbK078SpLg9N7uKgCKBkMzgrGt
oDWiyW53MqKA8TtFTAGNjwrmONkPQb0cEBpiPpyKfN+PuqhkOUAlzAYdOsLBbDaSBp1kxGm+3A/k
UWw8vSqnS3Qdfyrto59IXcp1/F9v79O2F/xf2DuNdHzPMpMdgK5fN1fG9SAquROW4zoFr1w9kvws
xRTj1j65QMOmC7eQpYq4ZL0Mx2KH1qHV8fL+LCDf+DbX/iekQAP92LP5Mtsez5N0aU3tBkAmG6Uv
tm45D2RNZ1T8W0luZrhUWVEMLhmUFJDku5ppKgbLgwsYUjo+saTtWnLUBQXolk3haxmS6F5Z9ACo
k9/2xWldcSdEqC8xN6n+oGgOpxSSA+OMmcCafLDCr5YDQwIiQvuwHt2Lkyp+kKz5WO9HE0xGhfTv
i6ZDZP/3EsIGLy1nl+Db0XvwtKG9JSvcaAk2P8PsvNgIUJoYtkgvnn7b9TFCZ28YVvqWsYXnK7H4
WeXiZqPkZfRJAgF/9cJs/uMQhMQJmHS+KOt+OPuN2tt2IOZrEHcsbQT/uC8PLr5hfOryPzVjJrRL
dyqzBccuJcKB6T72W0YFoLCFXNYYilOjrnSiAaV1XO2B5pXG/QhXzp9RJGs8N8AFTB2a8tJyzMSU
oEi/qXbB9sd3H8GGg3QRC4VYt/BicIne0SqR8oWI2RYTqPST3ryBbrpIffcOynApro66FUH449kI
M3pDi4kV7kSmX6DttQkCJSpQ2RPOtCA7KyiGk+9TUjyZfbV4xl+B6rzf90/v2dS4lGIqOWjHeQKu
BXZszMNBPjzkPqvIYQX6EW2fYcKGgZuJ7V/Pe/K89yxmiJQoSjK/tOLJljndm3/vKZoVvzdhTQkl
AN4XPlgs8fyKpqkc+fzfeGRiYWuDIKHXnLRVb/6iE+Y3p58zgTrxYkvt5PeV/OedvCpcd4jup0Q1
1etaXB/wdJxait1cnuunUo+pXow7hL9vjtEBKvN6jsPQxEDd6+rM0EA2AaoCyiNy3zd2viT7/X3u
4IGpNO3885cSehEZnQwbed84m//WgytV6wPBF99q8nEICz1fyrGJeUOqDRcfmlEz1L9pXm33yGLH
pEZsRyZSFxAvfnFZHX/SNFnXEmBGWiZjJ8Hm8icGQ/8Nwhg0xm0SUT1iiVSWoTbwLmc8hxf1AqmM
uL7OHRE/FBKEfiHk7L9YsE2ryrm6nvVhrxj0kEX9D9sjaGH3mxPm6qFQMKyyc2ozDBI6MTNgwhHn
4oBRblXj+mhEe6GNcfVlM2eGlRfPcLz2h7ZobiI+20Ja9U1v562nZiJZ67eSk8YeatMt5jPZmH0+
1CM0JdgIQwimqaS+08qe7pT4L7L5yAqaY5CeDJrtUBGIP43En+qdik8hyChca9JXcu8QN4EQ2ihA
IX0ucxzTXWcA66s8+IOx/5Ijo0lq0LRoikddNQFkL2oYLJafUyGiHTRefMk3z46keSQGvQygWO7M
j835Zit7M46xK9Fxqjll9FBqDVnmNpyzFulajh7V9MCeVIzHoEGjJO4jev82IrUsgCfG2U/BFwXQ
vZ0w5QmXWis/9o/CgrucvNNDWZh4U2P81ZTVSAbN6cGkQU222EwuKXs/lA0tHCn3boFJ4iM/ucHp
NMFZ27I9xzy+gNwxl35Nu/F9vL0bvgQpYtrNxHC/tSOawsHtm6tPh2zFWxX569vFRlRYTlNXp9gJ
3SJGvABHE8WzkECwSDUt7+rgBfh6FSexW+LEVwjV6t+1N5xNsOOvfXYxPw0Cn4+5A9xAz2gOVmsi
6oY1Cx+5G1x1ndK9LFXpBt2GlQAzVlJNMNflFLgVw+gr5uJvaFHVBPUwRdFkdfCvRPCSQfMIEm9g
Nv8B9Xqlxh9gME8PzmicXZ/51dYPgpY4SOlwIR6Fm1oacRBF5wx1LlSw+U4yiJf0rH/osJu/Y/B0
QTpWMCFGfnFs2Sm5JVwgf1/K4mUVgH+KyM+9TpCfnaB3assn/reW+Xb+q5x6RPARe5UQ8GfgqS9p
3CJ5hIAS7aq4FF1Izann3xdZ9MJyJ7LisAUvur1/6saveJlh1CxGKGpBF0u+JR+9TMPRWBCJggcv
B/UVDJ3CcaQ35fPDdg4tli+Oy8kplFxZq55rpkJcKPYnfNBzx5oQKHrDhPLNU4KxLrj8xX7Okypy
UPilCx9A9283UjR2RG8DGK3ZJmZ+PIfeJX1Fj+OpdEsZouILZTGAen4T4jflOWnEFbumgv8FoFfH
5ym3i6OhvOkT6jvj3IKStGATtyy3+9b4Nknobx9Wq4LDx7l0mh93r52f0Ui8Wd7GtwH/rvxCq8fe
TCh0ahISLJWyNWwkaI+2eQ3/hmbr0mgYoZtmDwUHPugPD++FJnCjhqyh1juTVXRieC9fSBdtB1As
YdiffX9NCeBuAgnGKkYLAVsQ0nkPCh6E0VOiWonnpfvw5EIButnmUHV1AoM9IzNMbaVkXy3g5gZl
XsN58PfygBtdPhG4U/g7SXWd/ENJw6T3lx5HpFNNFzIjIo1a8LKRVSBXPTHtDH7Kxr9TPAGfKEFY
5BDpAID4J/RoGS0UwZTxEeiIViCptv3MZJtazGYnsbZvWINygh5KJUkXCYPudxC6d2LiWlv4Tkhw
RzVdjK7vU4rLodW5ZHok3JhQ7qcRUHncRW5MjYgIhfMhmlVG6P/q6xTvmUR8n/JWcef1dywo1gmF
aBsUpUYi7FR+WgmZbDVUWyf7FJxVWjvcOl1J9qW/nZ4aYSL956woR2x952fyPEuPehZMW8/EJgTJ
GIgfj57agliNJd28vtJbt6ZBWki9Fj29nMB5cJbyOcEN39+Yv7l0LipFcynL3lpwEkFzhIswEoC7
O3PGhrwTmF06ryXAFw2AQdFmI5zmn8V39JRwS1PH/22aI7mbfQ/VMtkC4u0b6f/FSbyQqYTxB8eW
i69bz69C4gNpw43RqLSbkC0skFN0VjvikpBzrQa36PFWOwFiJIqULP7+fGz+giILUihA78CesAQ+
dynr2CTM1GMN9Z1nqT1ORkzutmAtnEmVjgeAeO0OPoEePPuMNqSdvqagvbiaySm0QDFklB3IqXXO
575wpFuDAfj1ofw4OSt069gGEs7ApHzR9oPtDm9/FPJHYLkHbNUeARxEHpu37tufGlVEPCPl7+i5
ekp8fMjVWJtABsaHeXE4NiXdzVX9iPU7ODIrNmfcOMqfYZHXA63Umd99neScf6psu+zf+zbrdGqm
EjBjPiiEjWrGhpFN02Q36zBJgtHqFHHrvhmx3jcEEC5TpLVOJ4sR3usYnM6MEwh5x2dqIy24jZCI
wGb2eu/xaoYRI0BrJckiiCC3L96O21h/dEqlrVw6NH46Rdt94XT93rCZU3DMJE9UzNjJ3KP5DCsC
3Bq55rkjYhrMP7UGGV/IW23DaQLgf/Pe9FlXSmivbY2MEGvOYBt2POK6lMHkohhOgOtMjZ/qupLy
FynTLYDFpcqL5PFFYapPdRzgmq9at4f3GMhaqy2kvAKLenwld06e64/bf5F4IL8z5EZwr3OPTYUV
KQyievfWttBYgnIhbfb46i1VLPJzWF7lfVrOcZW/VBiJAxbQS/axkgUr+9zuOMeaJLRwDnlipK8J
NpP9EDdLJSzivT5Y27FJfnUUrXxoVi8Vq57KrIEmJcjgIt1RpYmM05a8nIcQHAL/er4rAy+fKtt4
co9h80v6tcwfAYqxFqQgzamLGj6g6YaTWtVQLForFpMduoQvGbYKP+uUykhQmiUDxW+2QI0UJmAo
SZMvfE6QEMQi6+bgvogOMsQM5G9tT4dryV3pDoqHn8O17WQA81OhDg6Dv5Gp+xmu1pBTYDNYZMnI
lmmxcJ35xnx/8dlIR44qQ+TVFX7Kn+NUkqFY3jWfXQtwa9SX3C5fM+6l61fsfQ5ULJry8qs2zDFT
DY/zvLNYlv4iUGNrUfglzFznewXjJ2jfVrDr3OXAQbI3oI0+NcQUw35CFCJCb8MOEvaaQElnFqBQ
HL4qLnXPeDNfABiFTdKSVfjg8Cga5Prr8CI02AV2XvvcznmrUmoPbUXXMQip/X3xImCGOCpBq1wZ
O9XE8F9bD0aBQBOWMY+YYo9WbbHiTcRD8Ystj7kv8uZ1bWdBS+fbWDiV1Ygb14O9Ie0qlY+8u83I
kU5LuR28unj1t6fnc1x529R219CKeMz/17tCa/L9oktFq9stltP8eauRnTZGU10XtOF9zA32F2GN
md+NZ9HoSD3dET7qAo7NySd5Hm3SbBsGKFi0BzYXeGqKSxngmgWyQFGGM4ruLOZbtPDTi6LkF+nC
0AFRhdR9k1HftZgM+MmhMtjElXbCeISrgO3X9EHPevW+jSV5MiQrENpqp1iJVkrQJrVeHuwOw8rh
WTG+he6iveVUmPPw13yq6A+8cN7xtDDv54fdWe4t5gY1pX6mFbTVQjMEmOoVaYkdccIELb7lsrFO
aWbRkzVIjsUCpBM0suLOxL+/ul0v4DxF/lRZbsEtaOlAWC2z2xhcVVP/xqYOUh6AeeJ3ozQJ2lRJ
of8p/et8YRy6aOXeQHedjW9CmUl4lIAbMLUUXlZlkzhoEUyB33RmRdp2p0O740ZpFwVDbux5OnD1
Ju7gPq1aBOJ3Z9sEpg1VbqXd87sVXn40K/2Kaf5a40aHdoEplvLStwriiJSnJI8R0IcvfKE99EBU
iCxcmVlAWAUaQd5FqPJyij+p7HRfr/VQRIJv2ch5qIbn2dxFVoTnP8OV8JsbJtQMMdVH/MIOVw2k
fBBWGf+p2eujNhcoaFzQoU2epW+jLbPpgiDpViTpoqB8fe2LVuJI2s6WpXPvxHKfjGi4cmnzmoOZ
p+SUPqdgk9BMlGi8aXa+tXsbLfIchcEZzfMDHZwPCqUucvqsXt2y+OrBCqdCKg7R7l+YKhS7ARI2
ZqDOh5rOoVZggsdo1VsRmKoo/HZxTdUrnhGTDJG7Qc9pKJNUdP1uwJuxUF/aoSqdUOyYdH8lmwuX
U+hGtbDQRhgp29xj/4nZWQ239nhQk5gLSilxCtV97B5+9tRZ+9uBHw/ojaP9lXQQUKZvK75xgMIQ
tPIMinKitwwF/ZsgJxRfp1mDKD7ok+NDpGZmMwEpAfjD1GOBkKJndEwBTSUEAp1WuSTWg0kB1AxI
2jiqeMMSjh2fEj386mTO+C1cyrXdAKUP7hbDKmfM4ZJk/dvpNoyzHls+1/uSrq33owWn4Iybqrwc
q6OwyloYRxLnMt14+lwgvyHy5EUBCiIi1OBaFAW9RNSxJYUvzC9L/5AAm09jmWiZljq4jboi+GcP
fqdPmaWwdSU/kXRFPJZ2bjBQNsG8uVaWHLcUdwmZYXJuXFxi/0fdthy1Z4Ko1WMFjhtcWKIH2mkK
dcd2HopGxy1vuIsvoTGOIQw6bol/44foda2tzYj5JB21P7qgpKXDla5GuwzhkIZqGJYxYGO+8fHr
SOW4P2xOnuBFzuI2wHutdTIQmwLpDIonbapVe1C/jsOuEdGrWZY3NGg8ELVz8AL/FFJyKDVdkw6+
0vMjTsdxwYZZL/U0cBFsrFgjTyOs+U1tzjoXud1gzixuQ2NIfif2XQOJCYj813j0hKLzGpyosa8M
2dX4enP1Cp51m84j73JRuI2/tByh9fB+CdrCDAFcwnuLNjqi9GmVzoRjlgphivlzKaUZlhQktwIn
DQ7wX9VnhIq0WWxY1bCwvjqOBwQ8JczPPJirvKQ35ouvwNgoEbQTB+vLHLywVn8dow3Yhr7Y5wmT
ufRcYpXRKcRJ4U7ZjFKaWn6KXgBwCu+C6JGnD1zoRlukz16viGlw38Y+50JeHhPwoBT2u3dNjTOZ
lFqbK2cvy9IPNmwgq3u14Ylay2GMLZWZ0PgR223Eq3Rb+MqHY3WXanoW3HVIxbTM78P08xu0BVFb
003sBZ3mMR17vjC7AxYoBI9N9pItaPsX1f5VqU2WKLYpYmKBor2/RjY7155hjzvXgYUHk/zPJ2Go
gGFZzfDMA1cIzc0vn6s2xkRdDpTXX7t9DWZGFlzkYDKdPQuddV+hj4nsl3degyU+amyj9q/gFB0v
ncijhNRmb9O79qhKBDVqKLGACdtW9VDY/DudT5nmVPE4fWWa/+wR8RnoyCyTnaOJnDEHt/R/xfaq
XuGSyTAeyj6RcoHYFOmOCxILvQDUYjPG221GQYZKMl33+5aePRl1XogTCiQWdjmTfEHj2BQcMdKN
npwf6NuFk7oCEVQmkChFtLMHvGFb9VFcFNf3UsKx3PKWTXROcbJzcX9t5tVaOxIwNepPKym1CWaK
sB5T+2jBCCvcDPati7etBSHNaA54i6xNop1FBIUWjcbyaj00hrjuEDlHGrWnK5rq5HyYzmhhB0Dp
nin5/+r/o2rGcC/5Ljgl3cP4akuLGpCawphEDa/c2FG0VcNrN2PUOXiyKpxdrmqgK3/vBbg5t8Fx
B6O+1nLrtBwEQwLjIte1AxTW06awqp0YlW9ns4RfGpcYbAoRYfxu5a7NJwqJi0sQdLSVx6rF5lIq
23O9VbpyXTmqJxodPl2jLkodkaEBq2hGEGmG80ogsNzCd8Y5+Jwu+M1gNZSmQCgsOPX6lU8wRZ8C
zQwrtMwm85dbqXmOYHusvRQclIFed10P0VR6v5iMIv+lI9CZ0D8ji8dg2voqM1oSmKyBgxxYjwOV
GnvAXTRROoeTfa7tbZzHrqXOOvJ0sUNxY0yFLJgoWIHg2VHdPzs3z1NEPPoqcVAfcvHtzQqyhsUZ
IIgWaJmups0TPhTBCyoxg8zpviX0T/m5zDGvQQxjxPlt0cppUY6SZMaqe9NgAzjJHWxtdcRGsgEW
s2om1hn/sqghKVX6O16ajyF5D3oV4KcGsNRUZ8BNWQwOWEpcEbxGbW3ElJRjrGCFyl1zw6MgL/R1
lGBCLpZKgWKSu9H3mYIT+lXkNIG3e0sw3TxQIohR7fDYeZHZXPsD8El2+s5QxPoncbZy3387Nicy
oPkXrMPhLy9Rsp3o0sqFkdcrk+41CCJZhuAIM8ZTox36SRLqEeLxIUzOna0sPHkrIt+WbgT2kNAG
5Y+CsRHLknt/a7lm4IVxaCRZZD87JBqFrJrb7NOmm0FZS9s1qOailLM6eIrwHcXfW0ShXfWqn8TR
68eI0PR2drB0qS+dt1W/4Cok8o7Kyh/BwYfzDYld21QQflzVyoVpE/2wvPsSN9a7Yo7XdR/6vGfV
hy3VRujMhviPVoqFLYtaW9k71PqXWXILAPAxMlnorLi3DHuSSafkRmoJ1JdFyje0J7ORL+aVkmwm
hmaqec1NiXjrR+Y1Wk5taG8n7YV6s5rN0CmcJEWxj2nuZREGsmJlUsaRM1dDQAHtsmR9CUI/LzrJ
UWSnVdxvBtc2I7r6nxoMopOXp1BcSEZo+P8sqR6A2aAu/DVaNDzHjn95QSldpDA5DWBhIw0m1zbQ
POvV5zYaVwU3Wr/aQfePfRzchg5x4uPV5OJXoafxSjXkWAGCvfU0xQLTBEaY9oRR6mO9bHsV95AX
ltPB5BvVELZ8uqx8+VpFEgrIHSc+RYsaotniK8+iF+wskh+z4ubFIgGZEtkj8Zcw92lS9s/JA75z
DcF3Jq1+0f0CINX4pr6WLZk+IE91T+8YdAj3Z6L4DgW9irCFxDu2N4me0rRt0xWjsQU8gjwigZJ2
35rC0dXghyzMXB1YRJJuzGXlXgvLyVZAjhqKcG159J7vM2eRzZ+P3r0R9YwgUxX9sQTL71kuUivu
x57MlAZjOymPB8S6vFLaWnTmi3Qo/Ox13GnVGvqwx/FSKxkAypfywCfSVNtlrfMpFjtyGsLTM4zJ
rWWwfAEXGqRFRZcU5EZsn/JgKIsM0KYnisw7qx15G8egvh3PN0TTZEOOazSnNdpuHaTI5iXV2D0T
XI7mt3fn/DOg0UHlgV1YfZk6djwtUCLB1oY8nUTPl+TXF/k3YQiKfiVCAHVVAimvhoF2m0TvS3QP
S45QzR26kKFC6xQ7Cd+LnySyIkdQzz98beX8R2nTGX+esv7+KiLmB7Sz7eqdfpNSdlNsErdd5Tpa
qUgbXkD9OQG2Q3++QWoj9XKo+6IMXTnmPTt3JiBI/uDe35M9RlGTIUkj/yKcutBEFGWYe07ND+0E
I/rPMSveqig12Zk3P2P1MXVK7rrcZ75CAefFYX37EG3xl9ibRpWPLTWLjgYlrFbo7Kg4jtakrANB
rp7CMD7i6tU6T0m9zsF8Z6v04MF2MIGbB7cUGrt5eSReJisJpKtpVMO+qIG7dYeLNyg4VJMxuCth
SMaJ/oSXe2+14eev+MKL87lj8PxUfPNQTKB/kD58G/DAVBT1RbZxBW8lrroB4M+DZuWudKJgxnZn
mumxrw2ls3pDc1VN9I9jmOWidtGzK/zQCT1LXvI1NcNgk9TYfaXyL6ZHHpsMuWfts5p146hERkxB
VptSQJ1yeZbjHu0VzcybPuw8/II5apxVAMgYXZKJl3U7q43ianH4dPjjLOxSCuicMW4/QyfYPdVG
K0TNMAFWDvtBV4x7+TGPPqC52mhhAhkLouME0A/jcfy1DByTgcczKD01l4ig7617M5eJmxC9GTIs
yll0lNO+6CiVTHMTYS3AEeXkdNpnflrjyBppJYA8pYjwLDiWgcUeRoZpYcNWU1v45YYhQgosXSZz
PfGFn2iGf8Q8M5h9HhX2RodlMmCWl6BHvocAGfVJXVehfF4VVNUPHu9t6uatfsKDZ/0kehVetp+z
uTA26HHtAyF53BTA5PKFsrts9zvbhKD7yt6aKXp71Io/9uCErDuiZ59xLd20i5juEh44gBI9YZbG
0DOICX/re6pxPaRq5pp3qr5Hwur95BoWE8Epvu7nPxLxQYXFrdO63lSlKNxcludcmwst0bOqjjZR
r8DjAD7IWBJ9gidpH9l5hrMEGZpTRbffHyL11Y9gkBYPYUaVD36dxvzOHvhSt3IOJ5/qsq0wDUZi
eAHQLqyrDp0mGb/Aq7SkMNlAp237HcQyCiC+n1k+5P0VGG11UaHeBQTpj3F7hlMKCmA/Y/GvYsGe
hFHx0Dr7XZIt/AqvL6kYQPrIUvfY0ptEtDLB7CnfS8Tl9DlFggZUdCZdpMw7Niqte/5j0HTUbFDS
efmi/OsCAeUwH8lwVfj2QNgqsyhhGuKynNf3AS/G+MTrichXKwwcjOqmJzobgYVSTfN/1nEn7aKw
iUv9rtT2X9PMlf6r76bWRTHh5FBj7GUiTLZtV4Tbb5dpi7ZXzsrWeLz83VcQ4s3HDjhrulR0mMfZ
FqR+ek8CSozIVf62Uz31ES5o/Quu3AkK+iA51D0aMvjruNNLMyDWeHWvjl4gY0PxyzXQ+KRdiLwN
l88OtA14G/pOntBRX+9mTntGcJVnuVNzNPTfDNg1CDxDab++/zpa1idD7QlDL1hIEYoSiJdWy+2m
iO3wTK5QB8cG6laEwwSEHAhXjaD9u3zauklI1eEA5npgGUwcSGvC+4Rv3tKRaKHojqVIeTHNZeaF
lkhzdfYGOOUoDsuMPllUdTkfoucF9SPKAvptOxKCULO2nWXl/7mD1PwIGcCyfEPmG2aQeNKsMZKt
zVVzE9zqD5b5kAob/FFAGCT3CD8z0FLfoWpdLeCLHbgnqZRtyxpPeobInl41Uw8IGrm8NEadClBe
Q233w0Dkla+D59cLT55A/szHU1xV3payS/4PIuRYJ2XgfB9+rlaX73fh8eZ2M5FULGnNGkz5/DfW
tsKfz7y1zff5hnMIoDF0lryqBmYDk9vtH3tczABkf2NKKnObVcqSf16YS71hPknqbUy0qU+EgSUj
Tdyoh1AkgXdaLcQSx4KKvMykjHf6Z4Rgix6yPU6vFweGeU3HbsScSoBb+VThbBhYBwGsEQtOfcQp
i2lF4a918MtWZUo/nu4mvd+jTUxFEzk4PTSZqFI+mVFIg5A5xNMT6RSfPDnxncL3k1z35RyfyOoQ
TIz4zciSu+1HGgB3YdT/qktnI1hCdZwCnscOyeVrqU7yDZu9WxtiLPhLej8KXoL83X7MebeXAyYY
n725qYrTPWLVzjNcjIpUUUwZoT0XajjmEuXD7N4fzGZBp3qv6VlBcqb9rSJnVLQ2p0P78HXmttzK
5lCSjPrEisEM9N9fWEE1Bifk/FuQwm7TVLppzM1e01f/XCQdhURj/pPgtJ2uZzZRJbCbaxeCMmcv
WRo9HXFhMsnOxjXUPAiKFYa1ybELLbUe3ma7sb9nwTIAG3/u0WZePWYCxUDNdj2lTOpid+6UjNlM
/MwRsr+wf7NgdOS80IY7QtUpxnv3TkUsrWnxrL+Nedn8Es3YoGBoz7QhNlzILWnCB7UnkQ2g6kml
ckHB0/4rbnpK6774+C1hTMeNqxgewAq+2eDLXHopAc9ZAbW5XKPs27jzPAbZJqRTBnpVdM1iBi/K
/GUDBClj4tneL2smob5paou8nUW9aYlpagbzD+cKSr1o47kYSCphu9qscr8Zfn+MCCIm2gt4JdPv
hYaH6dhwcsSI9ENjIZAT264yZ0b1kgp4WS2efbsimz4e/T3JbQJgGLag24EQHO1Y3IAzwcfdqvdc
NfLt77u+Vj2RB9Xeq9xZxAISCuSTwkwTOqMxDFpl63anOwO9S6T7WBy613kHSVuNgmBfT1nHBwq0
kBROhGO0kiISsYfJiUePRFz1EaJzBfZd2ZQTVOtzRj6IIqu9wayrYnBDcldtFoBBg2e2W9F0nRRg
orqcm1hiPCWgLtbVZUkx/Ekvdkxt1hFCyDxECIqHCWnvbbs75sQC2UyoFm3c9Dr9fIrKo1mheOO3
lXU87uBnbYssSyGll93VPVDcSIOUGKqyJGOC3bqvOlXJO0TBT6RIniH1o635SSasMsU/KCR/0KFg
RjJmJiJb7R/fhlY5FgHW32NHZ1+z2TRttxHnuJUfhjECeuSgho4Udo/NtudT81IfW+cphbKuPIpT
FdjJcPijkg0TAzxJVVahX2rKu0KjbTHdSXQMB/2y9Jt7RbAb6NRlq0m9IxuHfAsR3OXR7rtIpvca
IYrH1jz/Aj0YWJwTenSEtpbVns+dyPhDGkUkwCFNgLmbQ3ch4TLMepwqlmPKKCMrM+Ql5JIbPH4i
7jEvfFbkdJdAk1fAW2BmcJCYOdicZ65pmKfSaJYQzMrYoIjBg+ChELCaI2OLxHeT6KBlJnH/FvgZ
rErHASpqP9P6goSRsO4MeQYGKYvu8Zz7THPG5kgR7Df2K5x4t1/iGp7de0i8qOjOw1bbKRZgYA2n
F9yRw7nI8no7Z0uSZ8UZZobemg79sQXWGCGPPPF3ivExw2HLdyMCfUSWLRsVfUCEM+T20VuRaKGR
S5uHFgM4cccsphw7VWq0VGPAcWAjaR2LH+NjZbDAAcxIp0A2fhyxPEqse1/+GE+/6dKfnoh36p+c
ftGGR5qkUO/vWx8YdDC0YPpSfxaq+jaFEYpDPNozlrY1yRB0yVpkWcM/DmKLPwP+87F+ZUCk0QD5
Hzo5WC0RaHQO7Qcxf1fQ/Yap8sp2RS/5NsJxHr4z2l3w3xKo4imUpge5HdlU35MjcQHLsAiv840F
T2UqQwCvFsRXZRjTlPXQEZFIzv42tymrjyVfVRsLAjl/vpetp39w6EsTZtu6RvKaJ5ZkP+nxJ0Nw
Aw3N4qyeyMMES/hKI1JAuAg6k9eOvnk20gosG69ZUYwKNffb429ieP18x0xtfnpCax766FZ6T64T
wAC4FecXyKfC/9z6km+4tjl4GYFMClQBlSSNTKTrpDm7uXnoMrYuJZxk8JRRAvJphk+HoUufHD7m
g4yAyGZcTUr7nIjCoeyekjALobOSkYDn/8WCts8QOKn4HoK7zweUVbvIU0F9Om3OzWg08f3xYTi0
e+NblHRBVWEZyS3/qEFR2C3RW5Dw7PP3n5F2H48WgsPPWXi8GuAtWzHuWRd/9OUGy6cdClkmeGJ+
FzOvAxA+iJBLviPS/Qv6Be8ig9E+6Y5YyF+RGF3l3yaiYW9Ex/tgZRO5XNaDRI0C3xtMIdLHqTts
moKh0HvQEuJheqeqwHRHCr+Uli8NjBIYlv9FMswdBLCP/G38Ap+8ABzLXh9zAu+jt9OZM0q049FH
YTyeakLNnPw6xaebkCDF+/NM8lQfl4Y90W2IhJLshdjif1GHmC8qMsc6enPZphjjHb0queyXdWQG
uHX1iGxR1MpQToIVSJGjJy7fWVUlcilkYklWl7TDsET2o1xjL2IHkUtUJVzV4PrDBly1x29GQrQw
QXC/i42WbvAbwdLhmpZ2lc/E8VLSXifosRVCsxhFPFQ1V/P5hMW9egkk7wKv+VV85l8MFZXRSjXy
v8JtR2IFNBu3iIrA8IR3xjKArOiDX7Z5VSWkbsjv7AVQv91aE5Ld9FM5j0Vu9e0g54S1QN00H+BU
99MdYk5/Ulf4jV7yrzevRjAisiViHYyYPGVe0n9FYqvtQXnravE5taNC3rpKslj/Vno0l7PqT+ga
3FSvD1civJBy1dekGf+oO/I7hlCUvKKMfx9ZKgwJrx+3VnqdlwWni9yTP+FhKE/TWmGGdORRqqs5
t/y8/Zxu9DPn1o0971We7TUaAvjnYzU5sFYGy9NzMVdCDgoqyQ1z5n7UOZkTV3DN4EoemSrw2oOm
MPx/wu2oulL5tHjounfxAwlFA+i5eblYAE0ZdTaewPF2AuLn7mb/b61xV6JxclS6/J2DysJa7A7M
y2FXsga0akxgwUnn/SFao6lPYkxQgLBpG79H2Z7xDtLu2d7de2nx/6fcjW7hbLJSwCE8ffeCHkSj
DNpZrDTkQmTy/SopkJLnlWLXw40xM9wZSRhbonQz/225zQSffTQgfoegQRJI1odGNeJd6RFOMADW
sR+e8qXFp8C4L47PkUHR0aY6OiBJDV/4H3qJi/Sjtzp7dWfv4U0LdQlnH1TCsV8xPUMzrO4Z5ejT
XBxtrRiBP4IBN8ifM03/HyYqhXPkIe5y4BGm0MU1R6J48tEYaQArARcugLZI9N+fiXCFtkMcYonS
0uFZ5QaY7EI6z4dVaJcvYhyWomLeSgVwt+/0hsaEjl4wzVWlcqxkOuyh43RCk/1qfZ6KKPIR9/U1
4ScVlFK1Bhc6wzjyBNI46Cb5lXcF9Z1hCZbCrL4vVCn+PxHxwJ5Wfrw/E0RTIp++Z0vakH/1JMDN
/sONZpf9h9/EPXsQ6/f8GzDm67lPUTnHgkPR3pJwlp4zhXTv2llkH8NFjZHbm3UkRAEFwRqKTLtT
aRjOWQDUFnLddYoOPaL9x45a1yXdlEyEe463VdT9fzT3prjrG54CPAFV0CjJ0g2k/9YgiN/IU6u4
13IZuhDuygQNeO7VdJdvJ2gAzQ2K3Fc98KFt20/wLeVWrpA6DXJ5UaWuh5qGdEwlohNSk7YMO66o
7YwlXtWqC4SH9ZLqBjmpLygYxI+4tI4m0Y+Go5MNDCmksZfnQYKCo7znjceuO7tXhXBbJHioFZ2O
mzbC4Xsc3UWIDMtXslHdFMnCQGYB8PJ+1OeSS5FABPfC5yMtscf5LZHt3gKSf7Mref6Hq9XvIIcl
QxvCRt51ta3MwSot6a4ig5hOE90wtbTEvCkKIi6uYqlsGd9/gmN15wlTxRVvSGjPIP/G/Uo0Ulr7
c+tWLC4znPf1A40RxCv+t72bO5EgtGAp7h/9KiMnwgsGp05TsnlLJAFOxted3FSQnPgH4VxY+Ijl
+6nvFz3Rr6A/wbXdeNkxj5ZVkzElC06M+BNyurG4TitvY1YINefqmwObJhV/Az0z9PyA8x07/mAv
FaNB5qmiqBVPRdSFCptcp7YcdHcqplHg9kbyK9wyvb4o9InQSdS9Bg2x41DFaHCSZg5oSmL8ePxY
IIFucDpzNQFzJq+u7sjLxTewmoYMIQaMKpBlw5Mq2nldM1KXVkdwpKChBpDA/NQrYQimPkIMlMqH
+3wHr9nfclyIuyBr8WhNF4WGhi1lPtbVWVseY2lux/H+VH29bXsj8nOXudQtclMThlRQYX9piCLp
vKoAWfiuUz1u/q6qe8Pd2HA39pMtqYf8hs01MYmGJCnayvk61PIXMDHCsU1LeoHYyEoqVI7YyOwF
NhSUwFHgt/TMHeVG3Enh6ZIaC5esu6YPLBU5yLasODPQuWF7aNq1FpOxO8pNG8xg02RR3m72TkKo
yxf+HZB6FDUoQScb0rIfvB8atdUS2vzeJQfTcM5Py7Px5bH7Cg1/svBtufYt+/XnAcKAkElPbYty
N0Fru+C/9TxA1/P9/XZEq7ohYZ9v6TeCHVOlRqB8yEN/STyHROMKEgFw0t9+veSgqsVkYGVOXMbf
JTuFSsZ8/2N3kVwIO6eNyJ0/9VHd0ikWpQIW4/GyzissZcMiDFH2MVKj3vosGSDiuwzsBZJNOkZB
3sL9TD0FmoMS6UByuSeaueWa3tBh6KULQRjXixyxhIEwMJYPi6A7veY808oMjQb0Cb2va5KNrS0C
wjkIERSQdSkuc/Jv+GbZRMmhJ7N1FuqorDXhmgAmlQZjO3Glp9tTcnAOeOqbfHFsug8zxIzE5n8y
GVs+G30uAyUuT+Ej3lj4aWv+iAb23dI3oTfDSszr/akAX9Y6S5vUYExDV9hvzxKW+qcBVsByraJK
9+2ICqpxjhRSW68fz/aZlxeoi6qGpK5SVERGdVQgR2dTqm+aPpdoYrow5iaZlh69SQq/lzHuPegz
eJhcvOd6tQzQ/4hvHtdc15in2nvxHm4pX8c7rxvP4+A7q1Vn22NTXzKXCkXWrdVUTQADzreV/Yfx
xcEhX+RY1D4MpqIwA1dSI2DJo1OjzgWcnJo5teLyN7663Wo9qXp/O7u0i6BA8ULz6dUXL/MGmqGR
NquRpD8irpP8+MBX+0YPXPgihdNDp1SXvv5IdF5akVIocNvn0YyhNmhtjPahchZj52cw2LE+Wr1A
/I/USvk35HldqE294I/zHzIMPGFQAtDslz8noq8r9qNMDh8G9jietaHQB2EuQg0IvOGO8xvBzDe3
nM//Oy6T0fvAb9J0FeL/CnTxsYp4xKCJcTyJFc7jEUianbJ65b+cg6Hf2I0dkezFtwDJQ8O2Li4k
VQ5/iMU+XEJU7eDRWn40S5gJPxhM+5r6QXOuGnZ4DoYlXhMPXp9kiG0x2TgasrtB2tyyMPt+aYV5
YuvDtpi0W4Mh2Pu2dL5Qo9o5tyCM40BT9cnvYfEEy+XvqPU6afCL4Tg97029hEtcTk155XCEBORH
/TTK+F/N5ObnW0X6hDY7m/sC/CWvLq7tKRCTOeO/0TkHC1XJKMkkikvNkQqDzPIk5BHZeunwhAKe
YMZLKag7Eelay1J43s1jkBFSn3uONAD6yt+SQCeGBWFEUfNAl5XtbE9epF4gMMM4WAclg7r9ldmD
Nyl67xQ187EL/YgFPEvRLg10x7GjlTj0JB7ihktlVROOsDCaMOpaxmRjlb/tx9l0mr4/bPHjFuba
frvloWVyNUYq1j3OFE78uwMnNv7Xhjr88mSmejciTswO6q+/uIU+lDilh1icorDpuPW72IUupzhd
VoUcsQpNI8cj+gsFwts36lHcusDz0joIK9557AvxpB1pDwKl/nFk0X4Elup6rb0KvpRHBVgduGMR
QegLTdGjy30TD5oteh9TymEpN1//Ol9+28r3id9JVz/RdjspiumST52OM5YmCZyIMr1Gw9PiuySJ
uFYeOa4aOym8tFYhkCvBlFrvK+HwRKe39tACRRg65skiHjRYW4RVa6AfKhL8AtWbN6IpatveWgDq
1XVglMT02SCzkg2ErQ36N8aR2jzksTwx8R3tJX07tvgn8u5QycgGVPgoRMsb/olRJvy+YVAc7ADS
4IlXGrvf/10i1IzsOpobxe4JxtCtMOEO2EfDRI6wBVsdUXlfJ0ejUKhyyJKgoVCYg2mJl1DXJRGx
vUmHEdOvJgIcYHaiRx3v3/ukP8UpqLuoTmPrTHt9wVWEL/8AQuRbAiUogjkc4llpRjgVZghVy+gE
8ULk5z2nqwTzV/yAVQUgQqMpQyFhJwcEW+cdVyLhmTB95cF2w1dRUAczhmci5Qo3Ucaw3zsclZOX
raX8wJIbq5aFPhQibAXzBWyAgamEvqIlp8MLNQt2BCUdW1wMwdiSAB/URb0sEo50NbPsg+AwFGDa
yJNMg5Vjd01eNemkufW98R7Ycbh82t+2KQ/VZ2+VVXEGrzdoIvNa/O546SRAEpBYLHK7ZCDXcwmS
80GDtrVRpj6vgNYHoJ01ENItASKCY3+gn66fK9KLbVG7ZMwqtD/n8TmQrb5EhkFumQ82FFgJZpTV
eASWIEk7f+JmfygDZqlZBGd6b5hkO9AF4iC04xIQlBl6euvkwsFSvdQ6bbuks5nwUzTcLBsNd03A
e1c3yfIgySrx/JXlcSjp8N4Vs06c6UXibb+vKNA+L348nE6I+7wHgCX6jX3QoX5hqval/N+z8KJc
Aeep+gM6FQ7NNIcN7s6hf+fB4QEWYgijCu5644mlQxC9a7gIyRAVvVXwvg4cd48QOIzgr5RZDx7H
5DNQ4ZPWk44slUCCSfOrUqgGt/zEtBGIdbPBfjP2oHpZDoS+7ks9MWJ5mapB/MdCXk02hCoG/WVz
LwrAtXxmTAi2bk5bsVeBU4dYoC2lwJgmnLa7OEf/qOp9IkV469MeYlyP7MydnvT01yR8H0ZD+0FR
wuK16iuEaZpbQ+awjM5aRg4O6SD7ReGzTmyrjndXLWYtwDV1YYyuqj3xE6HA1J+Rc2zRDdSnS7Cm
Ko31LhpexfX05wgOKd9akYyyl/D8Wub/RTfLLKWiNFs3oW5r7jZ3g+aUNHLAVA/Pj+TzXI5caP3c
IODwoePps4KF82YQKZzqKDTysopC7DANbikjR7A5oPZaAoaBgNC57bkeA03iaa1S9KSeS8W0xVGa
ng31mEUErKdel+cpBCmbduJzY+rCtW7KYWqM5uhM3WO9UXaqZafi462l0kNIQ6Shh4Zmj1k3i5qB
XV/p04xhQ7P5a8cdrgv6rUNkbB0TOHE1+yoKperIc8jllslAHFxS8Rwh5LkuhVYohTbinzOoX/OG
wJ8M48ZY8mTpuE4Ad8+iSR3aU8gtq26fxO/ur1ovbMY6/kyMq/EAxlqpSU+zQJZtQAT77UailrGO
y/NJdAeUaM4WJMbXOYj0v1m5iccpecHA+x6MoRt0mwHVQaYD8Gr3Vkl0Fu6Qg4+NV4sT/wJCpxfV
6HpqqujORnJ2fg3jzNhiKgMTYx52/fhykpSOXUwDHx6uCFwihNYp1uZkMRNxoXWExLRLPK1jvlP0
Gl9ndAa5gkgqf3gZ1prf5vWfUqq8BemHPVZJoY1x3JnCgOg0h05lrSVZ80fWroMuivepsfja0NcZ
gF7XgmEiUhxT4eCj1blcxyM7l8U3rmvzW0b1l7G8A811SKkUBAQE9Cbf+kqyT93KPzjBRufJJhwH
cBP6gu0WN/Fth0JBdxQA2JU2r2aY0chfT8O3ythiopYDknBV2NZlDAOM2g9jxa5ibyOQKNHLWJ2W
5AONnXnw5JVysCtWEUxbfBUCmOQl7fZpQDbH5SE7KB9VN8zKrjTav4Qii0JmaiXTf06o59IsFWpD
+WOMVIG2sTWP5gc571aQV95C2p3cpPrPbOYwaE2Rjcpl7YZmkj/+FBpfTc6yKLnpCfBTiZ7Tji6C
JMKAJmzVAx1+p6JOpf8ygtayJEYYgN+OTd3spV2M0BZczyjewUY6zfa/CZx8jztet5aRzEMM1T9q
KN8xzZNTmWl+c3/HPPXLjMG32nkytC5YNNfEU/JQs3Iohx+/8Cs8nrmCOlc3MTX931r42KPJPdf2
TUEsTnzCHIs2wibN8u7sMW0rUyH9q3Ay5WTO40ItiPjkMz6tWiqjFtHH6pdNMtHiBVkJ+jDMzXUd
91Pv3FwLGrbx8K3f4/LI5rM+Eb1Z0iRjBOKiAMbjKSLWhhpfVTOgqT40VvpbpQKZfW+SEVvJzl5J
Jj/Fln1N6aJTQFlpWyc+dcs2Yp9cBfcC2w+h8KMn5pLh+zEMnaLi1IVOISUTDg1NPG5vR2FN6LBj
7MYQnw5obYI3unICO7k9pwceq/F5sCSRkTwQYbJazLLy7kWOgqgWY0OAK5dR6wuQxyx8kCacrcgd
ivnzJ6ba6c/IcdYaDdR0gKs8vAUqloOav3u3DAwe16VZNKU427GzePxOqnf2DbQXywG5KNnd5a6p
r6m6GZzxX1Sv/w16G6k5pk/gVi35MxRqfHH/bb6TYpiuBQlt+9JprBh6TrT7I2Mki8g+0h59wApI
LzIsaczVHAdEN37C4puSkHa1fVmFAo0Sf3RIV3QkEM3iOkwbbfNRhFwfJ077mYqrsfH5+/qz9JqD
cXG2qyQBJbfix7m8aC89ad1mlIXJ+rNu0FHjymYkzPEubx//OK1oSPB8nsiDShnPbS50zfc+/xfS
BqN9L95NTc+hyYBpkur14tNlM/k+4WnGs6n0SAYpPeB4Pv1uWxJe5VxsPsJkvfivJbHekRdwZowZ
HFNOzIilOercjTvHCf9+cI25myzAzdZDGLYsseLWOtntgehmcxMnflZpHPGJuDfih/SmzlVa5OKq
NUs7v6CBLu0n3RW2SWXJY8TVCF5Z8kgTXgm/j3Xz+exsPy7H+nQM3cAGN8UC6fVjtiMfpV6qj5Ix
BwhoqPJe8bE38m1/YLaoTHR9ZLapJXuH9Ks3P7hwrzuEMTDsyuXvnhoBuazw3VjmB7wxkmCaabn2
tLgluJT2dmnF7VjEJ6YVHusJjUnM0gwfTQD+nYZA0DJEmr3Y5nu5iiMwodCeZ3yhIlIZmGuMjRsk
p4nCl4LNHaebR9TB8I6uxHaMvWjLAmBkrirMprNO//oUC/58F58ilHm3WNnph+yNlPhMQwGe4Zyf
6qO/tRrxpHFXPZNBd+iXDF9xUg4+kNYKFzJk6nqXGZ9iQWhGq9/7yi2WHW/cmKAL+loQ2+i8y9OF
E39x0I0jJpayFd6WZIyb1G8uJSCBqAsfh2B7gquUjvcRGG1/Rwx1H0mZH0Ds121WaUz6KYPKVv0h
ttL48qVHvvX2GomK4Kay+fRFZwOZs3GAUwrCDzIMuFdYYbwhHMy60BHoeQ9HA2KtFJQhSI5QsVTs
DP2OcnBKF5qQjFdWVelpQyMGgVrURjzSkLBCGrOwLCQB/X++pOP3Zmzr7XTQU6J+tV5k5YMASEUu
amqst7eaJEeMZC/BidoyW6vDJ65OAXXZUH0HjEyddLix4cZpku8Vas1GvQ16nNxaEYaRLZxPRbw8
JRvc0Is49PElyx75gWpQCR6Jjj2eFubq9EWAlSJxk5CTgY6uQdipnTGTmmSvJsvLs7O+UwwQcs9F
UOa0Cw/TW4zABzPuSkFgg+K3ig6IA1IoXaVl1u0Gil/9yE623H3YxIukILalAPuCK/xOJY/pfxpo
nQW8jjohQ5GmcGIwQP2n3V8xACIQi6IyTLxjBWIsRPwqiSGicHfkv3BKKMDLNnY+Ng7jUhO5/OUg
VxsxelrFO2YzcVUBII0sinBUcbKFU53Kcehm1xCWdkBrPSEDrb9PZDwoCc4rAKXSZLO6BKGDUtCr
9GAs8xcdDfMo1Lbw0nwXX9Cb94I2VMTiYt1M79LacHfaU0Icsds72B/sPQ87+WmR2My4CZpXsGLz
6bH1vUD2WVZ0B/DPj7utkqNGzYAYY72UlwjIg1XHM4GCQQ3dHcacGGxn27ugzOFmJQU6fukERCaU
/G8FzQm0iRTdhYTw/o7/KMk2BQUavxKfFjELVYPkFrR5Clft8i2AgN8qM2uDO22PplDCQREaDTmQ
4oCQFxrZI0WotHr1laUoVm/VxrjSmuo/Ul8hURGiL+2shl+3StG52FM+eFx2Sx4mlanFX0e5KIT8
9MCYZEeaYMqoT4CVcl2ncAjPwsupqcRq3nQ/2/Dgmg2WKryuyLepCcIE+s6z4yl5PYfx0bjIBEIG
YbsylpJIvtYN7xis7GLbak8MFognuHpCDRU/I/TM946ceTJqyby52lIW8z8ns5Dz5uRHOHKl4DgV
qUVIWy5odaZZNUvCP9KLvwOLnBBwLeqfFmJ2HPr0RFjOUXl+INTOQXrDLVROxv0Msz38+YSSbLo7
ZSrycRVl+FSgxRRpm01Sqg8qCr1X6lrxaXFdkV4ssTSNZDdnYuTz1MFAVSn2kvY8EOQ6C+n116Ui
8Nd+AgI+BufSmMCajL+7GgWb3K0TrlKtG0HJ+I74lDLDfAvxgAsGYcVIC3DxJSGeMkcAu4nYI89J
aJSMjuTvMrHEGf8j6gkX0rkon8XBv+zQZIrkdm82NL+wLDHneD++YnKLKGAb+UleurJkbqRo0a6S
HSnz0Mz4vvpyTW/oRF44tyKneFejrMkt+y9RkCgD0DL4aUXpv8rYm6p9gUKXRjuLIg3cngDAC64G
vMCWQ0iPwHZZnbSjABT0Z5o6DY+3lsV62Ujc3Vdkapztmym8TQU7BiRv5p4abhhP07Zhh7UB12mD
76afrp8JT4BhEHo1a3RBXbCSD2xc89FqId4Cc8ndmaqV3D/IVWueiSS7jnth7r56pUtUkaaejx0U
+sY2B/QCM1vBMwWWYd3EK7B8P31DVuc/q6hlVNsgMXmCejIDC8EhOvnb92M+M46B+SXvFgKK0sLz
uptbBeYbDefpKOyv1FO6w0itOceo9Btqa6LVsDzW/3u0ZbkwgBUwpcvScf0EsuM+SqXF8D6edcuA
LZ7IeNd6wF3lHu+HFPDDdsJ8z3Ro0b/83yqSDlwwzY9tkbPjf9fFisOrWnKHTwNqEVRSVsCsF5/b
X6/x8G/lAT45DXnDb9yJKi00+0AuVruW3JJerteDmB9MPp7Mpckzz7i4M8eEby3/t4benMtlwIQM
yKEwLqwWpIqYZrpMWo15JXUQR26u7/L56AeyTajO6d2mpfmae6F0dbHyVerrqnUyn8a8mD63rEYo
fHu1Wac7rvgvK0VaCleMLfXR2bKl9/7oK2NtaesaCR6XpHwJ+hBXTgKlgwdnd7SAVbNJpXmJZxP+
ST0zU4Y6FDpGoQ+R2noJtHQPmYMcxB+0QO4DcE1rRMsKBAad8AC0BiCDAx1Tt9nDfdTazZKnvXC2
oRazfJkBfogvNZ4q7B3xMsc5VI+CBFCZE6nY5YD1yLvFAdGvRLLCW/bZ/mp6mg7bzexXKiMnjuDr
cXzt1C4HG+xGFgXV9GQ7DF07vlnUCCrW3JoZ54ncqvxNuJlWaON3Fg+/hHUqyj32DWkpFhPKv5qG
39JgCk9rxOHfN/6SOX7KEFxO2NHraNPNC5uQa/rAAvlznm/xzzaEy2oDi/bpExrKbWQVph0zPHES
1HeHuJ9x/vwSTldiPIHvtpG8nXVqASM21Itho59vuUdHj56pgZb/02s3jM/O1GGCL/gSk+AM9gxP
qd2z0YeY7XUArta1tlHI0gcwZFZbCDeYGWuxgQ6/mjlXA61MlA/2VnDeic3mqswwrQbw7QMAQFSt
Al/H/sjEGlKe896wFVT6D91siEBF6Y+q2AtoPDm8cHWWOwJXKCAa9UBT99AntSA4KOF4VUefxUgk
sSdhnpueRah5osceOM/YMvvOUKJAkvAMc4d/hVVtC8pKoXk45irLJyZC2AxOMFlwsSnRaiNI4Ac7
/dMTWU25scE3Um5+QOgdj7GC+N1zXNmqhIBdnOGJo8JWH0if1ss1CD6KvoisVLlQWcjkx0D8gwwR
YJ7UdHzMB2/6pl1PfibSOjzMvN6FnVBw+yqfH4AXWhP3RbdVqPkYodkd1IP/v8roo+y2Mx0hiypF
UmZ3fUWPqrk3e6YVRMD1UAtcrO7HrlAv4QC+sVgGC2rvMz4M1vXplCOVIVNzSBDSX6Tm4Jf3NK/W
nKw2Hill5/NIWRNeZ1PhJiwT6AAX0PCGXwrHR5Sg2+iuc/PsGfu/Gf+l0VY28nfKXDJt2nJYu3Go
rrvQDFKbECacUfxZeilb96hADl7CcNCHgOqcfyIXELqDFbMr3awrelAA8/Wk4aknrPm/j8kogaEX
gXs7uWH8hVW1RHQUtO5an1lHZnJVpJtKv0UxNJHGK8M0L15uHgtXRZhGh/XOpJybVd9q3LlBXGz/
Zalub1LS5Nj+E6SkQiR0noyix1FzwO7IouLww6HNKBnKKF90RCdit8QI5yo6g02ZMrCYflPN2YDv
1Sx7DZfQt64L6CE5MEwFHTKpkg0WrPKvFXIZn3b3HRpAffSioaPiQMu8KwGBgfJOLmPAXMHmymYZ
rc5G8s8A9BK1I5C5mTJiKVro3o6ZWYC0FCKk7WLqme1NunCSHy/IsQ/Fawk+0n1v7Eq1rhL7G0wd
351vTYmYyGvRSzOWav8759ggYm6QAQzNcRcXMeef0wKTakkLczGlB2PUPVg97eRm2MrR9dx9S1+0
twstAIq101rBZpRamGnptlEphQN33SsloEMWJu+WKaJLUoyjWcrm53KgotcfSjA/jpJqIVAsdZLT
OF+E86uMRz5wNYu4rzX3ZISuXPMzp3IQHw9oLkn9aJzwOpvY9hqlHoX2LYutI4ayWvjry+hf3KJd
SVVu2MfJGw8FA/b74UOsBmn8V6ev6Jv48+k70wsl+ribHybb7n/ahMLmfSyVS0SnCiTIu5r8qIW1
+UzOgbZmjRLwxw37fCZ+5txBeg0ubjMF+RL+iZ+VnPhMvUqQ9OCUYuJ4U+0dCKPrlF4+bdXIz21s
6/SvizDmBAso4TedzF0aOIujZwES7xOWbWtqkshCFJk2IlCpZaF4aNXQrCRZnPXvVFHKRKAm9ONH
6oOMXXuMT1rT2oy8I7IeCSd1smd7hfpfffC7gMe01aJlZP67BuLXnkXcPQgVSiGfAiJmbVveRz75
pJ1cmpNzJj4fYj44hz96prJIyVYOLJh8qb/qQhfjFksIGLc76Lp3OTOZJok6+9WAU1b3pwlk0PVR
9DNbqvwSUrjfVJ33Md1yFsaXoh80S1z340tDnQTwTLaTSQEiRMRx48pbvu/Vx6be3/3Br15EOCW7
yp32XYyX8ASVEp+3w/T31bLosX/fJcPrjtY+z0rbsDHYhwlzQmeoA/NhYeGVZJLv4bIE7aWgwkgs
r0twGmc5KGJ5/y/IIunZLvK1MyuF6ZFdIOG5dHrSZou1fH04BchxJsPwECfM98PYb0pW2ORT4caW
Ml5EMahc25svuxDcdtf4cnt72q18uCO8hqslcm9n7vF9x+wOs4bEHV/yUqaPyLQrmzfHFiNRE9u7
sYiCu4hQ12OA/KPu7CtDSzPAxMjxCLjzcppMu5s5L0LUAc6T008BeZFXaZ7V2PazaIyEmp+ru9fR
WJdqV+FASznK5v7ncolow7ChWDOocfYJgM2EXunGEF+VhCsTm+AcNiy23ECO4nUMOjAzhwyQiu5E
QpG3fso+wyh0Xl3Z7OsdvxG+ISfnoaUPYFikD2MpkwJCLLr4TfOtkvmBLtMK33a1AatSJ5LESPhO
ZOO8tH9YdxPg2bBsDHLWW0tPzYPTZ8vxI3m2B4AVmxWTOxuDPWY4X/LP6TScZBRrdZXivju7DjK0
LuTb9xh61cJmwG3ktHIJJ/3L+8QalcxOP7SVuCeq5Qf/mUw0JrxAsI/fnCps6YgGKcRugA5bXjTl
J28HsdBE20eB2AzGqarZldg0RFEnatOh4GFBaTkJiqBuDXGHNZMNUQHQKWEpByeqeGjTLHl9iOY8
GJ8pDRWAmi00olrN9pcM9eNzGlm9gsIviaMouMVE6BuEhmyRfPzQohw1dL3IngarkGuqE3yp0mpy
pJpgf0mMgqxsAs2Gwk8SIk3KBQ8vff6c8wDNQubDinxk23CuAzeTw1bKgPAsrvb4DDEhvb+x92cq
QXAcR1u0MVIjxsf1R7Ei00ltl7JxbhaDuiAD1uq2c2F/55bUdf2AT8sibiSoLfNG91gP+A+w2tug
IZat90NI+KVt22XSyYQDZKRLRpQTP8fiuYRuLWKT2T/GOYCLG648FaLVcfKYmxknyqaLldUlxMVK
baEGCgQbyYyOs1FK1Qo6KrFDTh7aLpUUBnBvTnPilzQsiSJ08ueDO5R4tYruqqH7afe4lP3Kn70k
xeRkTfRjxlh8uAhPLcxTiPu6Smk3pvc/Qmwq57JRyA1VRJP5cMeuU234EUyVyYusL2PrDOyp/9ge
py2BRA83swfdsl999kr7sjaTnqyOQ2VyMlSrBFYYYi4O4fyu0Hnfb9w7ZJPojNXRPoK4RaUEzbsE
Mc95EWTLb+RhOJO2q6uQn9/ZD8aMm+NDlzn4p42t/YIGUXTXYJmaHU1ec6PAx+K8Xy6pUdRNsm7f
XcuyvRXvqu/DaUtAM/S0py7xrGFculAOELAgqYgLdLS0uA6U7vzyBNDESoPP5jzilSmTsxF2t+WE
bGopJtzlgyuTyHVPrtUQmyWu66pzi79PndBRc2FxsA9km0mTv7ZIXLaNsmIf+F/TFoHal0ZlGpk9
XlZn+8cC7YdFOERlzv2sEEc2+1D5ol9wvv87pHusJwbNBu37HxqBOr6afi2IfJn1COKTFfhqNalN
lqrYcnbDFE1FIpE7SXUVPJhnSwD3ucXbZnVgACAfH0uNEP0KQpLE8Aivamg0BSBSZlVI3uZ7OY6o
bXNb5PXrzpNqBDh5Yprf0a/9uMGePMZOFc8HPZT8ZDm+3eGDbvXHvPaehwyqC3aMZDweUnP6sRog
N8l24rfE12/VAd27qTS1A2gXd9GIFQCiWJu0MvkjUkzq6MYpFXZkMNyGkbvf0S9Hxj7GwbSIunVC
yZSiPCxsES/BjvTy8mI0OLd+3MURpU3oUYEqtcvsQAAke8eoVdd/solcpd/oBhNvJjufn5M8co/w
Xgti9XwJ+MBCX94t4I9bb5VxU9bUsQ3uvkudOecurweFJKyQY+maYuaXgb38xOU+PNKwMiRLLmHa
Q1PniVqsJyPPOzEVGr2tWvbMkK0qe+WvGbBBBwcnGtoDCP6PfESmLyNC+n8qlcFikEuugD0bDJnp
P6owKC/3GKR0GpTs/z6ayVKiqKkCKBqA5eapz7Mcv9BquC6yqiof5uPScnj7txQYgwbS7Fl2pxAL
+tC/s4bfDlsNKPiU396xyxi/tOMW1sIOK09nD9cFivDh0znPjdC5m9q9BtFqxkDX0QU2DksqcAW0
jRWSdA+k+CT/EEoXIYCpYvDFdHtifBRHr2aeAq2/umhc8V6eUFPjWfCNcV2iOf88FYHMP6L3Pfnh
JmQbdqOu037OfW8+rRwuBgLTImPCEEsYhmcK/PlJF5F+i9gKMlmSKegUJycJznbnUgcFU7gbdeaC
NXwGIcL7NkMsYuci/MDiiupSX4jADakIfbs5TeBGYxjOc07ebj96muYCMcJn58AVCofXU+ma/BYE
Bmn7AEOgcQ+x6yh++6QcspBf3cALlgdkkW3fyw6RYNiCgLez92Z47wxGtjKSgn74dhBtgAVDTr6r
QQgXmQZJ4vbI3vkIvg0NJUp39kUEmMC7EvUo3K2PSgUTEakrAJwhHSOXXMoGC0Vji5tyd/avWhMP
N4DeE+f5vCepLuGiagdZep+/i6QOO7UTvC035RHvA8QLD4JXAnDbg4mACBwn/b4gplnuRVDVGKaV
xUaaoCPfZhA4MzgzYtcTrQdVh/wQtFXByQTKqLLbt5eZw7hCRd712XCJ6PYe8fWx3YGPF6qfN/v+
Qu887AKboKOdw49ux3wcZaVgtSUu/boGMhWyjTZCfR0bvkUQRCMg00RVJ7sXnJhp+/Bn0aRV2FI1
T81gy2Gccw0lcKaKQk6k389VovfhIfWF7uVk9SnTvZ7Lk/i6HlbL1xXyryy5qmV/YIzbenBqbm4o
+QAlDgVlnhoExQIY2/4NegA32FC2H7UtpGEWL+hYrcWDi5wjev5bwMCvUoPRiF/7UURdLH46Q3iY
kThc43cQl0rrgmRahsAg2ZLrmN+IwzrIHyefgb8N7/0obigh2ULm6yV+6xdWHotqZGiahgtTaoTq
HpUOyLp/RmjG7KuYMmcO3ExbxS1DF7WMZHlXjiX9qN8/ebkrghvzP0ZqIp2CBE4X921V3096kYhM
C3Okp1QGvy2SGUzLRG4qiPlSR3hRFKtM6lO07iIoF+IHze1QNX+uRShfx1Ml4mc6+BUezh5rep/t
M958SnBO7q0vN0rRr2jpT6sQN9d2qYWYICqX9GElWoeUXTBwOXB88hSVzKRUtyaJ+ROnoE+UKAEi
fuUiHwSWjAIUCXpZCkOF1Ed0EZ67U/juxTjApzZeIviF+R6Bd+gQb6PeSrEAIx2rDJEOaLju3YaP
W/9oz7JJ3oR23IorQgPk2lOkpCMCPWq252DPg5PBUCioq6CU01lDJbnWCgDzcqPF5aymAKwMA7z7
NxMWKFxIgawBEEoj2sGo2jInnbRXZbWv2CR0bMsQBHGxWeLcmF4URwa0QYXwC44hFnJI+tm0WSFz
JbdS/sOjz9NC7VoRlmCggDRw0qcJwmq4o2iWYQMi2JZWlaaVNhqB8YZ/TXSqd1iLJSyTP4jwyAEB
LHvP5HxZWPb0s1AyhdjKsnxqnpmnXvA3kKg2JqKJzhsORcrGHUcGO19H7GfhMhgKkV2IEMR/p/MI
qCTQM7NWsUhTIE4vyNTz4b3T5o0Fedt7/5IkXi7bSv6LyjbVd3Ip2x01UU3/5Jlo1lYDW7TQFvqW
PEXaJZle7EVBsXOiaKyioJP49FUIp1+yJGKy2hURJnmXhQtlbEnejqNvaJRYyy7NcIkM/UbxXo1f
qkmZJ9ieKHOQJ8wwUL8BAjsJPe2IDYYAemWce8U2EHuoxHlBZnxcsk4cxWrmX20Y+ak5dZiMJtR4
cB5wqt12XrdUX3auoXlNHDGrFRMpLsSHswGFGE15zE1xX7KVpkaERnP7yepPfhkXYj0LrGFitiEY
BUNAwoxKZYQZLm/H9fdwDtAX2eGM7A5iAAHs59scLiJ7kNTCtQozfEDDyl4V2xPE45KwEtZCsqSO
LeGPtbZgiKDriaXxznDmQ5PWpmbpXHurzeTheAPeZuKRHUQ5CbpTWZ1KSU6BGvOolaJI49oMg9PN
iwRtLDrm4vio8ShKlsxB43i0PndstmFaiKgu4EfJHgr/sBUYZkwzq1AzDpd0UMhPiIk129DPXat6
GwUxA6mWxZB8tZhGB8qFPNSuvlTLGqci6fboEF3fYtxm7vn7lQ/0SMrnnx2XyT/9pZSq98D5usgV
fQTXVQJ84GvtwJOmoG0pkAV9SVHAQ6zfdIdhl7BWHgdy9rU3eKfnCsBbVaHDbDsUAHMCon5PLuTv
C3oONUPeVFo9oqh9JYw89/J8qYA2O8jg+/Ay+xJuusqACPQCYGqB3qaXjwLqyAHgFO7DyreG91sV
ebhNipVsSuZvxHTMtt+oigfMUK7Ef/q5nSD+mTUvBbgrwYJZAgKqINA0T4ilo+/u3ET7YcpYQjWB
HflzQ11Q6tOtBmZCJtVRXmigAU9ym5sHt+g/vxp73pVMj2LVk4sHD2osPp09+KQG2MsO6glLDbSS
vFVWgIXLOl458DreALzhNMPpKT9ug4eow4mzC93xH+urKy9poOHBw6yVc5L0O1pQKf4b0b9qdzXL
QdJ2gG/jrlXImjCWi0ELj7fw8ZJWwW3AvU2wTmut4jPstR4BjI6QCAeZqwGsihYN5QZvlfShhtaN
L7Gzzv4B1SD7EWd0FnpGI6knwkEKmoWC7MX8xfGqqNfmIwfmhIkSXoEZtRz2JJgs0Q54DbERxXVp
Yl9N0LOV1nKkEQBbuPiicUnQAnB+nFUqCqXdJ3wkczG7v44QlhBsEu0iWB7oZytV1f/v4bwyuSti
D6HI/810XY/gzjxbBk1Ife9hIGIeMHTNmXM05lulJZ3E5xe3bbVpSds2vScykCLRXqd2y4ybIpEg
edkFIg47yIuPi/rPrnyT9nnZKFHPoeaSq6wr8JNpsCsLs5VaDpQdCZVi8aje3P2C8OdTzX57EQYH
RVbtkgZhY3Z4UB6hGMcFjDwny8VOQYmVjunH6CIE4fdLGrUUR3+UiqmsTqPd/E3w4yl2ZMtge1I2
tllocdYxD22laYAp5tRH9DDVQLxE3kBIVJXsWuk4reDXsOcc1dJsha1nQEb4BOIJx0aHIGK87UeB
OJ+e5OuklWaDvZuje+M1bbMaIf5M1qkPWXanJdxYfXipnOKv40DrrTWIQoPl5FIgMVO4I+p3j84h
UyGiibdUExxWbeNxmqx/CniHVUZCiEYDjLiRSTlXlg9v3tqwXnydCUk6Y1CINPOwoVFbojogRsrK
Ep1BuM1DGj4VPmfRkm5C2vAnVfrihjKofnkt6S69G/yoRS14GOTqVgN1JVEUTlMZfs5gRi+FL/QQ
u9AaznUHTKNU/SThSaMVP0gXGamh3OgwliJRcm1h7w6uoUur3FRvMLqQMvex0bs3xjIOZv7NteEX
Zn8ANcWWusfgJRGTmZlmqer4zyZkF1/NyiYd3KbCmPWaxs2eSlQpDTZMQgVzEwnNMtv19+vq8J0W
xMABCspoceMyCnUIitEVyY4HUNi0Kw6/XWa3VZSGJBtH8eVBbLBwKcrY0y+4UAOFVRWDd2yi85m9
/pOtq8yRfwdOSOaJq3loU19wL8RgIqphMvUpDHt01qPoPLXRUfLObMJK1JgYcAXdwlPqEpKLpOrn
YxWdClqqDMIBTpEMLMntKKUBwjd2RydgDBaAVTM4WSdfXy1wUeegOtz66l/x1INHhSdPpCXrrUMl
/DM6lTm/LU7Nt6cdRwgeUcVptkodMIL7AEtOW7FjMpbxy9E96vny1r8xz9R/WOi/onsFijtqrHQU
jOz57bPqqqD2SsSWkf171dss2e1euawV9HYyGz1kcuxQhVcLDWIXHg29cZva/l39679GXTkTEUw7
mguZcUXojnUBV1r2eeNwuRXc72M41w8fe31YTiACE8tgaFVgoEEguo3vUHGBijUhD1Z551yf9QyM
ikuxvpEIGUYiCnGLV06O++VW5jeBzc/nlqiKMdq0LuPRqg7GmhYj9IuICiM6Jx7v/NHYoriWu1f6
43XZfTRVDU2XYif1IwXr5U7BRsH1HcVzt1YJqKthYNbB/wIBGms6pyAt8dkbamKS2cNsDQSk2zrk
De5raDrjnxE5C8IOEpawY/NynPzvYoLABDptjEZ0ZyfwTs871fYoeJckA+BLAELOJ+TLQPZlVEGZ
CduUyaNC2WH2Q8XMEfLffcU6kCUe65jYTuqS+jfoY0QfIqmtOQHBjJ8PIA7ZSQscwXwGn7j+W7Ol
NGF6Rs3zn9u773lTQFHPayuaIITtA2QxVKfbAdX/EqVzLXjuCHRZ2pbr+tP35tJ8HrBoVf//H9Bg
qSK8I/JGKECD9cfqAS3zVOScTHYHUsiA1FBQvo6816zxsl4OkM0iq8ARO7rTpp6p0dYBd+ev+/6i
+M5aC7rWAyjt38nTFT4LM5LH/2KjfIK9cGm2Lzxssh7iJjuWKDg0ZQqzHIR7b8T/zRJpXZ/uKAXk
7l3gGCtkh5J0ZnqUbXh5CfJmaPFTQhbPkHm5SPA+g+6UWFcXV4V04PMHHugY8cDyiPJXwbqx22po
qgeLu0+XcjjkYNSvSHFl5xNdrLLa59U3a7nJQVWRIY3PD++8uOW/lPDk4IMthpkLQN+h1sZqWXTA
aX1esMGxwdn/YEaF2EqF9P4Xs+W9XUzZOg2q9e8kOLbd3xfAhjrpRb0O1PbPNYPbyMiXTuGNDp9n
S2N3kgGTvRc4d1p5fdtuZ41M5CNyU5GLnMw3llrFraHkAlZzGIdNLiqFqU7jbtVUoTWNEnGax0Po
pHOvafOB2lfyMIzz7trKFLjKNMoF+TqaJ9koXZIe5uoJcDYsyqZVnV0rC4Z3jjkE6y+FAOoohUFF
ci2niiESlu8nx0+J1S4S7ovMM88x12g/JKuA9X2BtDD66wiPlpUvQjdbjRPI35hPQN/SG5B5bGap
VCOG+4vip2JBmjLi0IrHkOaJ6NkKMYg5VutU59Wf9DHRqJ25nKL+QPmA7vSydT5nWZ/0IkgjwEFm
FK1Oe71XPnKiks5gX92odKshp+mDXFBtX1QN195DOnL75YEtWXgmNxRaS1x9+GEz4xzjV0I1+k49
LvKrP1PSUNXacHQ3LxdPKU+LXEz5cvJNvwQIgGRI2uLI3bNPLRz6teNgqms4yo1SCXdKTLQUuKC8
rfy1k9Ccm27S5TaFRG531dLIOJK9g/VhqRLTGM70CZ0o39/Uef1COno7xJ71Bas8VvSI30KfAzb3
OznQpgx8z/pRjbbfR5GMPrzRmKvLDOwC2NI764qpflydpUYnOIMfze6fguXrsjG6SkwH2NDSCkrh
qTWykLQ4PsMISNbDuUP68/JtxAYH4pVuh2ozyPu5oS9aknU1hU+nJGyhZWHMS+cL0KPmgMwFfwBO
NTSoTBSoujxdkJJHzZCa6O02VceQvWWwxDy/mLwqPMmiil/vN6CdVlSofmVmqBTzMoGalSLvT63f
w0PAyEzyeYqkMjkhMB8etOq3Q3hbuKsZJ5CWLcMqC0mRxM2Br2rtemJ0Fb58I3ikng/RygTn32/e
XB+gYXf3jac0+tmRTPhAcEoEjjEz29XaBzFwPRIUQMIODygg5CYVwFISoJWG4nnWQaGcG3RiWGxV
TFCpVj559UALNa8KOARcM5UEQBuRI0d+AJVCHgCq4snAH8UIPtwA6i2K+lg/ivgVWhKbjf/GTfMM
SmHMtRzzZl4xkfxsfFw+jfWPxqEOjUKShcIBafsQGsNy4bzai+tbceKsVfBSH0buZb7YNgYvENaf
TUDUIJ1/2fCJPXyuxd94F++GzQyj/XTe5/WLrAQdi3hRovxPDPVW69SXCSlfKZxd8viILCkQh67/
Jd9XoQBc7AxD9iv4GQE3c4nmbBTOaTrm9zT10+zqACKkqRhKbUSuAtLRgAnsstRztB3XXunEFtwZ
mm3+6ac/Ln/otnBaFL6KyTr9xAIYw99HfktTtM+MD2QX9YXC0lsuq0JK0zakU2eg0SXi+d9WGdUH
RVTuDPUbZ7A2zRjgE8Q4wdaA1bSWJFfmpw3ItVwCqx4MGFroPJHpFV0V8FacscacjTaXEnuySZ8q
JSO6wr49Qu484AyhdLw2x2J6VfVyLzcWSIZkAz2ayWbLLUhQujev45oEI6wzxQsizwdFclUVDSIi
V/NgOithC5C0sKSUHtj0s19Gab+zKNBjCTUJpzBFnVq5MucX3gYWLvmxB7g26IQ3dp7nmAt3B/wV
6NNLeKPvIAD2i8c54RC/P5kpVoiiL69NdTG6H1xaiK7a3UJKVA8I5gl4Q+g9wxOdL+UVDfdT7Eo7
W6lalXdtZbZ6a5MMvNz1OXnTo9JouUCaiv6CfnZevZXr5VUHQqdAI3wyR9rNU82fZ99bB/K6biFc
ENnvLB+w9u2SCWKQ/dTcqFEX/1q+mgW4e49TESP2VERh3JgmOBTS9syCG8yuxz25BAiP375BJGjX
i9z1o4O4xYHD1rQAhYttXFWTbYJ4UeCH4VUh+327CcIxg4+NI53MXODDIKXW4bYmIVtcIdiyiDpD
AJdbFH8/pHmIuZmpU4fREfxRgjLJQRbfOeoa/XCMkpqBB4Zg68VMrKQGTF/ve7zwOat7N5j6ShW9
3r02NDf7631E5ak4DLeaRDtqMhiFjBrk0DDGq3uI7aYRShBxKpvLLCBa7xOuheCA+YRosz+qf6+a
Zg+xY/EKq9U7vCsgc9w4RgLvre/djokYiFpXa8u8RwuYGS2HN89w4sOuH8R9AuR2vUyckZb+UPx7
yRiwWhf/G/e8OycZJmkx+ej0Mqpxf8nraiv1CcF3LQCNcgMJiyxIhiEntA78YlYAWZanCpJMeF6G
9hxg6w+uO8d6b2ZixNKCy4U2OMdDil1KcVN5k5DO0+jRgZqSN0iRXuAbJuOn5+6G4xoM2wR+JpnA
lX2F4ISv0RFCKtXwpwSkcslg3aBcEUct8aIXZ5xQAeE4m1WLAYkQoFEYKqjMIBXWNALKA+M4f9Tx
hPz9nvlzqrTQl+OrZrK0QEfmpRjmcve/sOebqtQbkiK1rv76JE9lqVIfxtVq0nPoDaSxmabShS8f
6WVLsV5Jk0AgJh4pR2Z1klh6ue5bSM0Mr9IaarpI5ecYSXcCXHvRvWAZ5UvT/U03J7dpdnJXOmZS
go30GTk9UUrvn5RQCPuMXCyVa9uYZM9f52csSPAa+hgoq5nGssmXjfmN3FTszGvD6mEPiPd3TMXT
MSz9ow2eq7hkoNq3aoNwOOgREWOcx/S3XDFDJ8heU3sSHM+rmXCGz0oGfG4RvqpDGwzpGJlFnoXp
5ZJYSpEmP7dSAteUUma1djkaTVa44z5W9KvTTK0im0cuMrSV3T3vyOPWyjBsd6cNZdDbFm9K6yx5
SmWyuBawsMgepQEyb9G5c3E6Cn6HJ4V5WJ4LE2TLqCbqNHUG7/CIBy2N3h/rWMXg3PI8m/mx8ayx
WgZlxIZuv+lrm3KeeHHM8Vl5rCXoLS4OeeXRrCK5N9+aFI2NpznjdBmVjMTC4HOKToPPrzoTjEI6
nLnJJoXhd8UUlAj5EQqN61WCPpTTmkUu34ssBNaY485SDi6IKssAS3wZX7JD03AEsgcYoHGpnC7d
Hr2FGjw1RSk5FMMbNz10AkTKub/NIzAPnguc7HxYm3B7MKtsaitCnVPN49Txqgy3JRy8i1LB+VW2
ww7BLL6VUBHtzpgV2Z651DQ5ikBDiydHTyXZXr0Fs6OjAL6S11QSg/fj8I1ywBhlywtmF8wIPW88
cjHbrgMzo+ozDt8HasFF8XM2Sz565hsFO+v08XldeOiM73kURI//aNlVOHkFvIcBOHwcJHhBekq4
vPYnRrpXYBL6pcwNQUiA9UkgS/8RHw3vzeNwCSrZH/aW7Hyiq/uLqkbgoX6D2TydFjMZ7DAti49f
DuGBON7G/9It+iENV5bG6PGVVpoXXk8dRhs2NvJaqmXSuH3QKc3QoxUPN7Unp92Zim17vMof7kxP
PgqIOc7auvO9HyOHCX768dHK1DGwtf2bNrFiXWIKBMjGWTZREtw6Ztw3aPymQvVC/w8Ywx6fBDsB
/hy+mDUsV/tOdSmyD9b2SFmfGzQs2ebDihQI+hoUtE12sgR5kt8ZjWDH032IkcsvrZqIuoODUBYQ
xi/8leCtg9jEeNLGls9ML83ngxe5IgqCyM7lYur6i45HpnGK3VM6dk+iiCZef5viLFSIZ427RWr4
6/LGhvKtGXGNDHsWX5fJOBq9B2SvenCkBXF0k1e6Wbz5tPfijsFwRVkGHYzI141ICfDGMq5SZn6j
aq2u9rJKxV2OlxgXGDMhfvts6XgyBzkZKbI6mxznlHFyAaiHFa/Fsguo08RfI93sjVIfOtQkEAV/
rjd/2XT/6kf99bS6Jx6SnKDhqDKQ7zShHmQhcOQ1+bd4bEuQkpqlAdxmUl/HClQUoRw6jndOtuhi
bL/B/cXxENEoES1P48qPKuix8xYqKGVKZ1CEQXl1rTYvaglc104pK4e2iY8tmoq/3TjjVpACKATu
9JFGSpusqR6O4aHmg3GBca5O4orAlPRmN3dqKXv+6JqGK5EYLehtqUGTQt33AS2EYpbI54Tgxd01
Yy6C8kzXYpAfKAvFCQh0j+WqLbCR4GMRe5q04wFbxfSJNbxBUoSrZN5bDZAv67Q/PIPf5V1iL8g6
j99/lE/uDNoIkjwpsGy7bwfJgibYKs2mFHh+Jdhe3l7CvD6SNh43i214ljot9G7v0gXRwfQNw1ZM
9+kSYI0S1gkck6r2ubgjagf3Ks969tsnLTT+e1kF43PEwsvtNkvpDfaQAvwgFDB1WBqsA+9nCSHs
tHq06wFM2T4pVZb3vLORC6zu32K2yTDlDdSHS7JiaA1823ZTu4ZWDvJu5j2Ur+zFUV5URfQ19yUu
rWjzfy65tsr4uZmhdZ72fz1EWes5bGwLu1BseiF/9GpUWdSeAOAe5wRCaE9NzlofYH3T9vNZYoUO
OzkaGms5cbpmAjaH18lWQjrYK2MFZ+HxNk1qsrZRQ3YLegPRAGpE0BRqv5BephnXf5FViRaBSyRn
UD+meuhqHstAMS7WUoA6XHJbuy/LnFStvyk0jlr/Ohy7QJ3PZTH+DSQHrbke9uZJpJUDasz+FV9t
fx/JpNlyO11E/LXWLBl/9O8Lpbp+fS3acCxpTdXuAFRjR7eXuRtNaU00xtpSW1DhmrPxVx1LRw8v
IdwUnMlT0K46/czDoGIqru6NQ9ISJqqG7nMxlXysIGwFy1iTEu58T3W8FggbByIcG6SvnMFZ79Fl
M8HhtJ/4GBNfnBLuGTdTL3NlQPCuKvK9Ipvjx1sgzX/0dzBtEPXPlX0QnsYqKYuT86Pwnm4UIVVh
oMGjTteMsDBEz8CQLOf5zwK7+3h9YV+yZJz996X257wk27INTgYRo2f9n7uNN2/GUmbEVAfG1yET
gsrjdBHsFC3bNFaO4ENHLYzaFfIirnk1t5z5gzwVMJkFbiJCMq29GDWGy2LAuFsTuI5FBdPX0hqD
KipAXDROupPVoOBCG2HznxGTbN9dx1y+DcHxncWC/AONgXMS7dXqVIl1qAgktDhNKkpeNT+GT8lk
ilgeSgJzIt2ow3IHKeThvttTzlF9Ac+8S7T4uprrRJ94wmxb3dm978mz0zokaOGqjqgVAYL/G3EF
WQUyg0RfLpN9SwUqAUv7ZoPd5NTQDOkG8sVYOOn7yl45v1RMgXk7aniXyvT3ds/kc6XpQO6/vuVf
Nz2fyw68F2zLpJxfekOR0ZvI/eTddsS+YuxiMnTxG8ML19w9Duh4OnlE6hK5YVQrVtS04Q9/vZNX
Te7YTKxS+lKMverzaZ322qc3VXAWu1qEqjjTtZPxAV24WT4bLhneTHvehB3ROJbtxOuRns/Ia6aD
UkzToHBYcfrPp2FubikjSpuGwMrnp5LkLCneIUjZsTtllID4hFL+89n1WliFJRUqEJVKxy/4ujB9
ynd8Xywlc3fgIN9EflZcgo+EZv8wEJxi3gzcK3C4OyNilTDY8ojAiOb71+yf9927e3P5w8MZNmRO
hhvP9EDIErGAgqmHEXVcaskntHkq44iNUIu4ITcX+WUfOADkxc0ihroyT2HfG3QHea+eg94h1+dL
McC3DscNQELpT5OyeMs0x2hdyLMTEGrnA0VibzfTS7BwZPCE8aCLzfElvawQGjegPf9GwyAlmTD+
b0/QTuphGhDKJMT6HAcgJO1cm9aKrYlfEbEC4vTUT8lHMRL3jiLkkJD49TOJt23kVRaGKSmx+THg
gKwzTLYFPVjMfYZSoHqOkGFaHAuDX8NRVeoHDp9vrJHmBWzZ0HCrToR1ZTXqXFT9Sqb2YI9Bntim
GXnQuyqI2f91sWDCLIOgt8i0ueyewjIsWi5M0b3VHll/5ucFwogQRJWTQHrJkjI3zf6nCMhrR8zw
zurTQ1XvTUUH/OqmvuTouUnRzsbaCGh4KdIfHqOsUCLc/UwfArp2XIRZZhM4si0DUpSdBOth9jXa
GN0sow2j/S1ov4plW4N1nBFoKzt2WtP4KJa+Suj31akVmKVt5J0ycSRrHqZ699JAxGy8GHncKI0I
zOehQNAPQ8iwcbbY/zwK6OU5sjqWkwluSoxTZY7YxjH8VYtvRXBA89cpGSdI9Yxx5l19hyocL4tp
LIzg18GH5X9A5aL/KPAJoiaU29jXAuAcOQ1q81qYm6QrzUAi+MIgsuOQLAKBX9ERH1D4DIxjH5W9
H9fqFX3Xqd1ARb4yJfHnKArwo+1pVIcQYsqD1eso7o2puaVI5EKZryF41cNRoKi7Wb+cAVgSkeWE
/0Noirv/+99bXwUv5IICIUVNbRDaNF/jkJjkmuiiJi5TXs8GrL/0dhjiewqlZ68vDilE4Quwh5FY
CiRtrfqiwWkUmrz1Pjd7w1ui34mHLfWZHeB9nuqSB6q5QyiYoM9uyRzHSUckuNljuUa0nC2sfK/Y
WAAFm4Hw9TI1TnBcgtfCLfTMahsxIXwXVCmHZJZu01luhpnEtfCGklqGEyqaz8j/f62ACC8T5+SZ
jsKCCt2JPHbG//3bxmxVzt/0WfAcgBz1e/KTaagMXZXqoGG4djU7gg2iDA98YimdSCWm0KZSo3aU
f7PJ1LgIXfvP7y15nW/r4EeI6O0KLzdr9zMcXLQ6jREi1xoIW2lTM6qV4pHEKtgufc5SfCfVa3VC
Q4ZuC+S++e/5tgmO19DJh7FlnCE5aiJrPNlbf8NiExczt3fS+F5lmgPLmCG3DLeFUGIiZqUlj6Md
h9UkSElQt0LHGyVkiXRGD59xKs71CGZ64w590pet792BIejFDnfBwhnnZk3NO5+BGqvHbiuAr2IA
FP1P/dpTlfQe/OI8eCsBGeR39yr25GgnVCGlCAkH4qI8PvFjlU4gbqmpWk1v6++ari6vBzXGwAIg
lYjVY+qbh8Qj0oY+bsDtTrcpKtZjmm1u9Ql9az0q92uz/BIJx0yNUGNfRJIh0Nzj6vfVSDFVv+0g
kFyvEycDcM6C+KSJZjl82a/Tb8bH6YuQ3rDW2JOsV4OayYkMu8mSdOWb/y6Iw46Vji6Jr6UccT7V
LQRfoYg6jzXbWdXTYJucBFNzi/oCmY0QA9MKbFOe9wRJYl37eVdN37OPNtl8EBfYsB7WPCTsemLD
HwAOk6NlohIhBkXlbwi8GofaocRE395yDmD95dPBbZ6nxpyYlSrI4xZMC1jBGOMDkP4CQjst1Ry5
mzKNJ4gT+yy0/v7a9lVWtRnSzAOx4NOiadVKC8mWu+Yb0ItLl1ikzFYsgWPlc0+Ndkq+Utr+TGak
RvwKPn0c/06W6yeT4S3g1TRMD/Rg+7d/rdQp+68xten+lbf/+xg9ZrAyUXIns9IBip/8c6dTCa54
9WPxWgcSW8C2/5jWH+r04cQDh1reiCpTLB9LGog7b87zrZuen9F9Z+8yoqsxmrUTNDwFs4t3hE3F
C4dU2neN3OJTrzU++ohjDMnxQHX/hywUJYabusKfZVmmM5WW6VYZwnU07DQdAKoM7gZvwQNM7nLp
Wr20/QsKjvyZJZyqfPoX0pj/dpBj6WJ99jfm1hMjrUiklskU0O1I/PNssa0EvXx4PRYRQcDDPpvy
cOqQukWwfA12lOD+VWm4fpnz2f9FlmhxYEAHC4px1PX7xEig6ICmc+91oQZpqhatmFT1ddO6NFmy
lVDEZz3s3soYE15Kxh2LmcJqWn16gzgdLg9LgcJNZ2eaSyWcG9YNgM9w+3Rsv8rAqJN9atJ/XtWx
mVxzn/rbxLT9DI0eZ4qV/ydjmyfBuc4nDeerH8sSqq7k+BNKnNQsZjSJ6dCxhxO3EtE40pWR/0re
aXzLHLI4qsePH1a9VwrHTtdkkrxug51hoJboTFxWEY6Cil5rRG/9KtsEQZE0jKc+HJywggGCYkU/
4biOFJZdP0Str3JjpmBXIJ28qf4Udb39bP/HY9crxXdN8vW78/619eEXo00t64I6tPoplSe8mbXb
KoW8HImBK/btq3Zs4MUMboB0Qx1r2aHzG6vZNUIaM2CFT7ApQFEM3JqJgtQs5/az7fxrCT0SQ5yb
cMxQ+2re2HJMZh9ChKQ9TbdFwTyyWYw1siZKgXShj8KnNfA/l92OL8z0jBwzYEBdLjde63n8WEMz
8lOyV23e6qarjiT1ZXok4c0S6EOqZw7I1pM+UGXNONNS0FoYltxIPO/gqf7K15pcyDVni2v0V/iH
ec+bzkWKHJcG9z7JFrSDh598nFU+TQX17KUzDhjy7XG+kwy34TO4cC6PCy1REyWx1R1aLC2PfVxU
ZzHe9PqrK2QCQcm3MR/bFNs+ln6wODvWRr2iSbSBt/xbBOg9et35xxhzJQz2lO8O6/F2TxgKC7ge
wVZwvdXtIOawi4i6Rt3aW3CtghRK3rk/JtbztpVzBVhVMrRo1G6NrwjdP3lm+qgir/VaeSS7SAt1
KVvJzwpEi68A2EFAV0yNNk6LOVqyD4dAWQzXHUhSzImWQRHsEXu0C6ZheuGVKfHpaXXHKT6wfX4i
pC8SNbK7CJyNBJowAEigVpdBD7NT4yErhpiosmyYTXn6+NquSmY8lxHJirtry7D1PuqR1CLP310J
ZoOZnDhsrS5DLiP8xNrral4BlaD/yN5RJjc12DC2uVIdncifc8Lf76HvJfAIlK8BiDyAP71Jx1bc
xQwsHHagXpip9WI4afouKqOgaJ61SYwKdBsb/HbCFwrdcjEcMd1mfsyssSo4T+6yYMvSbA9zph1g
kAHwnAq0pH6C2lnkAYrfzOhCDpKC61RkWmyxLpXJjTbVLOC3mrjEtOZBNBa/u+TrfdETmJTKYGf+
rQzhSLoik2hh1kDAss+VKtwnCQSmSCPD0ZeVmmCwDDAN73AME5lULhH0C4b5mGwUp/D2XgT9lpFi
fDFZjj7B+rxTkTo0X2lakZnm7xS39KMVnfbzsmlRUnSq1SCm/+x2qUmlvYmduZDO8KjYX7E32e3j
0ewc1xG2NMLMmMwY6OaVYe98o+jTh6J08q2B84+1JhGxBjNB7plzPpYHryr+hI/9U0lbpCJe6Op8
yvwjwmjsYOoNNsIvjHKDemHT+yiZy65f8obFZdeTeb3/uEGFJ8ZfbbsW7AYQQIKQsQUJyHJJJhjE
UfAzynZlxjlyjAOaO8oix9JVV2fELRRR7fUgHtjQ8LnoUwVU90wD3EI0SdNrzLMNDOYvxDLsRGni
KG7wILZNFhcRwegh3LUIuteW6zIxZRoI3ugET/dh+vPi/RyN+oMq9+pwg3sutG4MlV/XKeh/FtJT
qADbWxHBC/3WWt1VSt3xcsF/24sXVZ+rcmhtiXQHSEUZoXbysWjwLgCWuVhSIyfbYU2ZYQyRB0SM
39UDG6PGu381/p6iuRelu6Y5QyuZHWaTV14RbpzbgeMQZ1U2c8pxlCwcJPcmwJXic+sCnVNCc2nF
b5FmxzgnRAfRReK3jsMREmMmCiyk4cDnEYPejGCvisXwmTlYbZautjvhTTCBJGKnXxu/WUL9DE3P
0DobLFE4dxqUudEBTaegzSjZ+7Yx935zEJFckXlOovzlFQBH8fFx3WojhHFTF2win88dqxo/cR9g
Y7AY3tGbTjW0y84ezsUyvoIsNsfARIaoQdBK2PKIBjl79HsXl4KLHsajig8Zv4WLpibYKENyx4K6
XAorAKIKHFGUG7t1yfurlq9MoPmWi0uEjX8td8iOD3+zf11KiTv5Yg0HL1yqkiHC/5x8hpBvNgcx
337SAszuwAUsLkeTKpJE1Cjbe1WyBwJjjZTjNER0WBnCqPRi4i5NkTWiHuwwfFJqvipPonlHlSJu
jGAsBN+XQNQ3LSroxZlkpr4flVV5gsseflwhv7AOl99NTaHfZFMfgGajfmxQmvMDpYwbv6oAc9fo
+5fKd4U3hxThLW1C7Zb+r/m0mizy4kp5pjwIXHGcbmw1c6/cFvmFlV8z8Fd2Dt/ff0WY9ZNYuGYW
zS0pzfpQgK82dfCJspXjFVcooM+siK0OVCeGe4c0dau3sW0Xn2T6vwcE3jIgnSucP1z5L/8aWe0k
HT+r4xK4Tzp3LPCC7uNLyko2gY05v4Cj+iNUchmh4nUMsaDT7Z1x86HB2kR+55AzUXbnRZiL1xVr
02aV2Nn/aLnaCpOVoSuHme2qnPGurF4lnJrshQocFg1SNxq0zmQxZxtkQ4cTEs+QjMuglV3IZo2d
J6umqh8BbN2zR7i4NFvRbNwE7/5MZ15moEl2Sk1LMDx+x/j4l6Vu+diVkA/SFX8yAtU/3Z8y4V1O
YB36cDumGnJV2nsO4O2zRiZElBhMm7JSIN6XG+KB8uw+f4dKgHK2faSHKT0ngxKLMZZelaANOwX2
wiT5dfPBVaXcZic61sY1b1m0dZZALa0VfMyHVPS+Xctse5bBrS+prKuWJy0wvf6Qcogtr7ubq2uM
C8mxdmZWGI5JqqfZXYNQHttjwCdepL7Sm/0lF1/ZBd00RK1MN71lPJC+JsS5pkxN+5sl1Vvgc6s2
C76eLK9k94VOz3I2uq5zkB4ngGOPyFaFT69FZVE8D+S6/ZNwvEhNUvlTrkSYRmeRq4lJLby4bvav
gtiGleJ0euqtPkRkJkSvWvcFm8p98e9veGYIXwk4kMOE00jJzIq/Zt1D/ZaCu6Pp/UsE7AvqCWPx
DgkBPhmQXYC2Cefy8JMU+U7UTMnDCoJwocQn52CD95Qm0MLDeMZI8y/YfwESYIm56kuhC9u90wmh
jjt7yc4Z024kuLL3+rmjMheGcMdVqu72WxBbKIQRgLcs1eT9Sep2/9ahaVRLGDnbV5OtZzSUNfj5
o1Sx72bEVVZHCuya0HyZ7pBnRGbPW8erZCGuJeZURXt1iPKjNxEddeAhVDTm/HanmPnCXr36Q2jz
PHKvlGlQmz9j1N449DF82sMwbqeCPfBhAKuq0fU+H6WBOSD2mszVzCpiOm5kCkILfdJ7I5EwMyos
5GuA7WtC080MHT8aFNPz7wU5pKeg67koPgF2Nq84AqSEKr4j9PL77dFMyKzCUjyVGKYR5DlZNF2l
OzejuhXutdQljUujJ6hDa80BK31y0ErYuBaD8yjazMIiOsPkjigotmjIeOMC/LJaLyxW8t/oT9mz
JWOwGXdlbHzxtqYIY4t6o1SGaZX3MrVjn6uUKzvJzeNso342WU716Ht9fPBMV4Isu1XIIjJ25g6B
31CousT8U6tPuPOHlXDjNNtEXGiaJsvyJvNjXxMYKid8NoPRPE4StjDRzm2y3d6ttI3P/+Rzy3Ix
4w3F6WSySTb6NKmsm4AAnwSgR6naqaKInoO4knXPczSgQ5tMNW3TmusMOo1TGI7cSyVKcun/pb9F
lJl5u9fryRF6aDzUmZgZ3BUYrmEvkj0LA51OU7IfAWFS2nhkit/lduhlL9XTtpPLeaMmNRXCWwr4
RxrH49fSfQWUimCNq3sgiBlRm/eG5Jic/U9JDxBCC/xAkf7LG1ZTNpwLU09QUYR3tqN9WqhRwHQZ
Pcrwe7S0JI7nOqHgfpNyPVmmBIS/j8KHfpT2tMjcVqO+ElUTswUlov6pn07/ZpTbmF3q96QTMPR2
6LYEawLChtY+WxPRh9WH2gXVFPkEzQOlpRmG5J7E+vVO+TI+DvNenk4BjY+MGUkHWAUUbibOecy1
bIM8U5LBfAxJkvZZ8jy0WKwsewI9+xV2XMDZ/KxT7O1gJ3pFifMjl5USt0GBQDrvgXlKFkXnc1gM
XKRoxMujdeem+apZePYbbELfdxgaq4Yn2QTbwk+V1I224LHWMyt9iz7MQ2oeWydeHcYGfxvwnDmZ
uYj4ul39s6h1cPRHVQUOA4mMbfpTBNf1lSexd0J72oB6btWbUGtRJlXNtxX3phg9QNoiwaEx3F0D
foBC7hjp/ezQ4xVqUvASeYiwatinJW+1k4wplBKUAXHMFliFKpMpf6ACNisefyZ1eLXzEqezbgA9
TYb9pZY+l/HxRSYkJT7TvA8qIv+5ONVUvH7T6vZ0LonhugKB70swW5m3DFg8UKekbgxyuCH4wMrS
HZMAm7MhBU9gvM4zu83x2yyIDrlxWwjkIzd6xm+nTV2RBtKYv+FhVPtTh83ioo06CQ3RAepQlK5j
yTuAb/esAiZGIEasHBuTqT7iCIwzT6ZfAE1B67WK91xz2FXrPqHRa6IAJOubE7AT4h3MHc0sNvVP
BP0SNBdHAPPA0vEGYC+V+XtpmTN3aIX7jsz2yKcuarxr2+MhApHlnyO+k5YS8LFVFMy9Ab6ZplUW
AiZsk5gX3dWBgfVNMAexZ3ow0zkCmc77dKwzRkbq2VgXjANbCRJgGfsr1NCMQlO5pQcRbw9LqDRD
MgLoiuiVCg1pT6FZD0QL6E823Bjt8wPnb+mAE3bjPMAkkBYUNFU288bk2twZZYHw/HrYGalZthYf
7EeDRnIqVHh7FJdG2/KQUr2ctXXej9bJsuhBXM9imFYSnbEVUkFVhUGH91sMpdM+3QwnOLwA/wwb
I8Ey0Ky6FYdEGjWYkfGQG2gEGLr3PKPmK3z/kfJ41WmOurE5dAxlN3bul2FobjqZbTQUCPn8TJq5
BVb/nh4DTbgg+OgH3X8FnHoxUFqYeS9uh70AZ0ZvHzkZFwXaPr1xN0J3qjSZATAgyNEj+q5UJBea
SKJ/3cPESNdHHUXAz7jzAAxw7pSOHIaImv+njZrNKyISaKx/ds+7xf4EhS0OfB6R/plM00VFXrXQ
WPrJxbyJpYnqQgzezIB3igs5W+CazEMmnuwJR1HRWDTcfJkoFTcZi+xtn1hNewEoGgf+nLmxFC/h
pr/KCuyD/nsxPd2xvY/iAooMSUggL8AAj4Uzk/WukUEwvyvQA2rAWRaqq4mwsXPTQ7osVqd5KvA1
gxXrO+qKCLk2pw0k+yIbGqK+8sX++NVGnhmELZMAr1ly07uO8lwEgT2P3nxttMNGcSUXjq5uOBcc
h3eRgG619Z7s44oPqQgFzG3SGVJ1nX1CZqFSsI84VfNvK1+FcCXoeKpfkdqMspHMZHVkpmjDgjTB
Nz+/FBl08Vi21KmiFTqkS4vahlSrXUk/nq2rUFECdgO1OeAtu3gLKkHozd59f9w4GnfBSZzATzxi
Umk+PbgBJSjxpeZMJtzJDdC9Xq/qjWdWwqy/GAGJgyvPzH1t58TYqF9p5YxomVnyR1GVYmOD0P39
RASToMn9K4jfyD2hxiOZbcLA/Vkjddew520dHndMmkbWkuuqsur5LFoGUmU/157whG0+UybW5X7n
rh6GCQOJ3RG5QKJyz9GblHzc7v9mFz1aYOYgqS2lTyYcrH+pWKs86+VRw6yzvLIcC4sIAVpY1XMZ
eH/uAP2A838qoBPl+v1bFbBE11k2p8eE5Fl9+sa/xQ2H9//dX4KH+sVSTocNXJOZX0sU55sN/Lly
DH5zQc+GIvOrFJ2mnaphAnsarH6DPNU30HW/6FwxMjZkzB8T5K1VrOO2v80lNo8m9MWeVrXsjn/J
I3IOqPdEhTw8IrNY/6yFyF3NtxACoVz8AG/S0WnDeVqyYE4iR1AtL+pXqvvYZeu4laCOKiIAxn7i
KsS5bYBrhftHpXffPP2t63ic0jhPxamn3bJjsYWSMKareBZKjwVt5R63zxW+qc7MEVsqvXT8aJ+V
X5yQblP/63oVJNdTC6CDCPvGpmfti1H+9HcjwgL73UaTw2y1cNMc0KL3RDICFuYwYppyaeiGFa37
V0hw/WvR3HXaX/khlvbOo8M7HAJdG9cspm0FgExJOfk6LmIi6baY1Z91+4p1GraSvnotguY/d+kc
+gR8YQOFJb8yUG9E0yt0BOOMft5f1e9AzW5hlHHUN7d4GWJsKWbRl8RadjHAU1bS0LU96pCv/qbH
vfQR+Ayb5TL5E24CbexbaF9MaQR9mRRxdVebHAe0NxB5vvsb7WIqNKSZAl0l+CHYmlVjibg410Ro
LdrnAjRjw42H0uquWM/nMdqMnDTiCjsOmj1+B1iBswaHZtvxTCawrcM1eln2CysRjQ4x2pDUvjpI
k0UOPAPHEDxGh5cTUk7qnzP9ERILDg9UbxSAkqPflfDk3+cTeMW4ujNpINk52dINEvUfpPwttGD2
Yc8yw57lgoydYtDYMoQVq2Zde1L3kqNYNi4xy0oZeAmD3KJIDjbQoLh5yOojN5F1U1mlL940aGvD
Cf9BgBhqj2q1NUSCmCgjnPYq/Z/QFdXhRxlMGCU1bMUrV0p17AfkigunACEgJqB5zcOEvC7CiSAs
W2aUOzzoT9Fk+sHVvKOVEm+e1RleHbrueLCiJ6hNVyxqmMnuJuJz6LXyrBX78TDrA+2N22REz2io
tYZOWRJUiZh9x/IZCCSY3IFH/BENPo6osB9742zLnzuFVgZIB98zg4mqRHK3M8pNuApx3X+Zn4Xb
BkB6ewOd0wosq4qAuleOuwuLArP5l4z8g2XSmsWSUrYDYEyz6wqSlfuVGYtCO3dfuPTpDSL+FQY7
m8BiTqRYV7vq9gvRThxQ5hszcGkBVmCkqaKYddRXY9kdu/0fRKpEvIC0yh52X0G7QE2z7cDfuj/1
aXi6uZkUJY2zAOG1Ce0hm+mweneDrBkrSfHqR6CglUxXIx7+RqtMjbqIlqEy8/08/6k6r1Dt23AC
RQmX+xT2h6euZoFMJbbjTgKqnDNbyebLSk+GmBXtoaHravRRl8xYXz35FnJrKXCPD5FZyEXwUeEt
vAac8SHUwyUTdT0RVV1TedWn2F88J4+xVq35nHSoXtik3BhJxBbcjyLsRfyOBRFauQ3AaKdwR2MP
84s/ZhezPxHhpvsul6A4ixr3GBQESXVGWBQbfbW+OpIuqUkCGv+R4tDKXN1mFSa+yieOuB5A3t6z
T/vZA4TBDaLqij6uuslIKWKrnwdLbS7I3oCWH16NMNM000e9TkGDhyJqkwpI3THbbfSN3PX7H/PE
kiVrXQtM+GGpgGR0D+Ans5xHTfdNewddVJjIsZ4XMlws1XXESFCtHIqaF6hqJXJ8OqKYwEPN5O5K
O0+oPhcOJyMRW0ZuOnVKoPrLDjYob9Sr9sbjbrcZzs98y89zKBa77a8U/uYLoSoQJ7tf50XTOepB
g8XPBew2RbL4D02JNrQU16scT6Pr1r81cbU9jzW9ldO+AkaQ0PcShMNS9h9aVtlyKIRmNk6Igqhm
pO/Ao6ELXT81/v5YMseMNPxo4fQRE+DuPL8OlC+JoReHbJDlDbSolyILy6kd5X/iecpd5MzFVewG
0JdtYFns6N8D2FNQWEKfhaNL+F+KbuKTj94uwsZaPgK2Z3aacGj1VPmbg+k5+qP7siZb/izsmNdG
Py3MklBTL9e1H6vE6BQcOcJMQkaCJ6D6kHb3Zim8LvBKNA0DnWt0R7WPWYzaLJBFmQDpnY0nwk0U
MWTClVkgzs2GH3Ugrp0fVUae5tqr/zdhcc01UZF6gdqCCWWEVNDBTmk5QTxKszP+Jx3UW5k48UmU
IYMn+C9U7xg4UgZvXwgnjhtwRAt9GsGlUOxszsjGJdM7B/39EuqQRhTRYtgTdiCdfedG42L8Yw6z
WKjuCFWuYROkWaP7smiEv75ymrKWbeDx/wudKxKNY7l4KUSAeVyr7r7stOvghpepilNnVhypO/HL
k73A6M06KaDfzjQhAxefYaouFPyL0HA2nvRckXLZod1feRgntIRRRlFCckItnFyB+RzsQD/WbaWb
SpeVsEIaHsyF1iFdi7mJ2McR4KSyEfopWlz51Z3f/78bJkUuvPEvLa0n7YD4B2dZ7y8Vk5eINrwB
s+QH3+Xbn46P+S4GykvhFIgDEQb3Go5zVOh+UjNRuVWx0ue6T5yqGH24K+YoWP3qidVzwF7jR0ob
3YiJVjnw8Sky7juFK2rMYsbS+Y92ccgzDuvl4r7+zI8CZd93LUS+lBV2PRVmvQs38WFHKpwTfQsy
HN/Lbm2fMDSbGFX68lY32P615WsPs/SYKO4R5Zd6iB5Nun9/Iog8N7OYVsxd8JlYNUbVmnTFELBU
E0p/+w5siKwEcv+Yughp8YVwj9Br48eDHIWxA/a1NICjuJH6nqyxwnn5OTwIWl5eC2+hUAzFYic+
mPYDd5bZKfVx1afVpS4KDyFSTU221vhUBN7nzbIE871kSM+E5Wi1sQQnq4L+fdDNBCtahz6Vqm2X
e3XfSUix+19p0cT1UBvo0AXyOkc/YUub/cJu40WP9HU5H2UrH7NmdcHRsRX0K4237RnSlRlylkmd
X1Kz+mlRTfqvIwegWur8TpTSyyDnf0j60bU/YOn4fL3XlZnS1aHvgpL6Uafz0z5418xHBB0zfNGm
RO89zZCdg7Zs4HPKpDG5F+bIOfJONBVHmZ9zBfVKvVYrIRTVPP0UWSJZQM1FoZtqSvujfYLrzkVa
mkVZS+JnXHpwc6vELWjdhpD8VaPiyEERKZf8tOcbY8rd36TeoBqqWvLYw/aSFyquRxm7vCZy2dC7
8h19y+CFPj/0nxlJeOEMl5m7jB7JT5dw1/iznI1q7NIpQ92kIMrk2NvCmFuZkkL2QaoxF2MbTNq3
rSc3e4SeUrWuhOpxB2juc7ite5L3ZMALMi5aNOKUOi1KgteYph4u1PdIoLlzzi7eRkH9lcRliIgx
r7GgsZndXmt0Yg17bCC5u8uSzckaKBjenUM01YOT4mAfq5YcsBB5Ox1tof5sxAyCsusKcyYW0QMf
QOYYzaTFUR3iLU1ZsN1WdT+QpWWIPDPNPXnQRJyyugp11x2U0k+AKXkkrsTZp6qFBMSXp4J1o+UL
OWaWF47KhE7VGljVQRgw/W59nhsmCDsH2l5wcIkvvgdE38TcCG4YIIieL3RZ1QkWjW6gqYq7mFCU
kcBSL2FIPz9A5cb63v6B7OsEqtt9nhXi6ZYc3WT+MzvFdTh6Ikwn3OTVxoSPaFunDrdP+BA019+T
/oStL2LqmoOJvjIyv9tL6OhH8c/rgcN8H0Pdr+TW58utYyqneZ3C1XDjnUtO0PBcec/9YCyeMgEw
YMQZsCZevDZVbbfKvdNsHP6cB7qWD2RqqU/9wihWL/qbhIGxKo2kb0FlSijGHx9g0Cr3CjCJe7H5
hWd5bwiezf3WNO52cAyOfRro3XEa4whcymg1UA19/rYqY0DbEGJvOlcdrjPbFZpSUx7RuKTVFQdg
kcxmo4BhU2qONXBJqpf0C7MOxkwM9fp0DxIL8qVEMPnEKLHa61NdTDzrdRRm8LiNdyksrmSfgSjo
YnWnVaeNGAlUo5MoVm00TnnWeGIl21azzpwEhyD1SnIBmEcm5CyqPaLXtFN294qPp7L1Z2jap3Ft
trbgjpUib4RHWWW31p7R7SPAI6Nti0m99ir29Ik3vKXt4aIt/wWIPsAsgYaPDoSq41L5eP5BFGKZ
0/xJTBvoPE20YWP92HKj+5AgCFV9u2ZQp6EYMYx8locftIyV9mahRAf7EOFd98pF/2MoIpAkcfr3
CxM1qDqrccq2myYMOoL7hUX+8RHkY7kIJeBLwEoffUCre5kguGKhbOC1WJbcM8sIpX1iEy9xcfLY
wiZ3+nniyH0JKcA+5X6s8V5WCmI6HEmwgy2jKtBCk0H9LntbEQ9xKjFC+ogqLptXsTij2xEEhtDO
SiGz2b6MeOk5gjWlyFK+rJ2NvHMz6snG3G6OM5Gfh/apyxEx4kg3m3YwVlg1tfaUghHPXxSHo536
8QV2nbfLpd0cyDKeJyOMst5z773DpEKJ5WjroasxE2AvPbNCGOpMpLQ1WRrMrEcGBpOLAerQnuON
/TeQNYfwGA2MDrzHB5RqcgpF0jD6c2vHSNBuW1qWIwxcM51UJkHw5H3hBfxV25da6kl2DSxKTsvM
s4Yn0wVYlRIJQSshQ4eLSgmkQdJbeDKG0fwDWBFeore2RyGeMJ+oMCevzUvcLpkMXjIt5FrQwYuG
PMM8jKkBBNvySvI6b0cXnITxn8DJp+tupCdH2oUjJNYULjRKK7tFcroq82arxh1luZgNyUPIbkeL
76pP5TQwAXbHCBVQqz5f3RyXdIbjZbhql8JOo1FBH5CTioNG+xI80GRu/TZbZjfUEUUlWJU2g/RB
e2m3JpCZveSOoTFk20xJd3QZ5WfHau+lhwtwpQA8pvjQsV8A60OB6X8pyUtAwYoRZEdvWLg6rwiy
FFZxa4SM5r/J9Qg+WEE+I66BG47yQ5wzpv898nnKiK+z1oKXnOAKvYBeGqjjxc+EZs99La958/id
s9wcrNHzIemUxGOjorN0vjoxYysT7dLfeXpuEyBhMG/9DqxpbQNoMeRjrWEdUCo1IkaVpdpKfqcC
PCgxb7VbiN3eRGWhFjpBiEPI3tYZ6K7E3W8jFezilW1NS7WJ5XLjRpHLj+j9skVtkvFyjdCWIWii
8VdZ3N5swVkwHGPr85tQkHhpQRJOi+DM6Yp4f2eBv518l1Joq8kAzQ28SeyGe4TdV1KGzhNVUjnB
MxzcWHNO4SQEk7mZwPta3ex65FWnLVUAXS1GJanw3P+sXkyUEqztnrqqO+xEkStyoOGcVcQNzqv0
D1PGvezQgxLAmXj02nreW8uXKg99164PyEjjzcrfWvClcssVV0p3ZbjovB3b+aFliKOoE+pOEV4h
0iDGsiIziwkZwsbwFQRyXsGuz3VuQChxmsztUs/TYEwd5rCwHyWo30lennO3cvt6AtZ5/B0jFlxV
CVwdwSNEZkRoKData4kZWxDANtB4iM3c8MI7g6yxbElaa2n2KPG9Y8STFGl2iP0x3eHXwmvDtX+4
MiR7U0pR3Y+PU2jMkYQ8hsPyyFQIXgNUKBo5JYi0MqBeBLDhsaI8wf0TrCMH/Fvcb1/QTDlfl7Xk
Ew1ZPmjXe04rPuJcnLFo1TuKJnGrfl04GO5MPA8i/a2MP4t2EdrmdRkSHTbNKDFXlgcrmw3XaMez
//zNDPllcVBEenz+STx05/CUqSzr9dVL779gK/R0nK+0xqTiwZglzPs15f5npBd2n/3woF+5KNW8
wOyKcyDGpf99cxb7B3cTvGgPN1pmrYr8tFE9HDpxiydnTdI0RyP0oRUxVtB+FdIIAuVhpx33N1dA
l0TJgZwJS2zMSPFn1yorju8rTmTxjU2F6E3oVU1C/L2f+/d4ZbPdOfe4cVWF2MvnPYee5vqedlCq
zlP6GRxxU9E32P2LpekLbmxBhEM5zBK9WoOadf9/O9CXXOzCNySKxPua69TAa+267GO+8RXyv7/z
zy0mJJM4UrniV7IX4RNPPNlgG04ndmdvqkQ/CErtuqShafOVUW3Ze5IAOgcqS2hKRta6RuspdrRx
eKXu9yJVB53mZCkIkao2D+u19tjbtoRgVcbINPQ22P0AYHgo7osLbQXq2nFZhHGgaC+jkPSrKvfj
K4TtwaUR9rVBmCjlE8hX2fgkWh71KXST8+H9rnIwsGxm4SO7Po6Vd4IyQ5r67Gi2NyNSaMaOdJve
WJRQP/TvRX0XWnv7iS6OvGrlXYVhWyTQn4XmWCqPjtyaRz7XzDCDJyny/BgZkwfEM3sywNHSR9w4
zQ945NoCdld/lEgB3SwUsFa+Xwe0dLsj6H5JtCdhE1O96Q5hwWvNuhsYaqsaeKu3QGjJuIvk8yL6
vurFxrww+1g3I0UMKgI+oo/PJUW6rGH21MZBG28tX+283/vLxHp7MR1dH274wOWRYCrIpxxZEtBX
TvmLGMXZnKaaEkVSkNFr98W80aO7q/aRqnKR8texfdl6AbtcWDXWfdV2ZExA3AxlicrKOc0QKfZ9
/yCnLF4uXxAMUPzYiGyRLOhTvG6JGAReqbNfE4nUKbI9UBFrJY6gtiZkJ/D4I8zljNNJ7pekC6Z5
FBQaEJFUdkOcwXB2bN4/GebBdixSxD3Xd17pzl/JY1eVlcgtjv80+D1JQ5JBzDUdD17UaZvcT3mz
orlBW3W2iq7VzsKdgKM/ZWkB+NAS8r3LXdjTgEf7yYnVMmvqZn+B4SWgKpX7mx01kp/T3477mGjU
V10EPmRuRqFUaHn6KwudI3hy40zsF8+TJjVmjJcif+9yOxcgjWZ3kqEzjEsMAh+lY/pQvVRbE+Y5
Hq8xJyCrsGXfsMiesBYStuUdGDkeY56WmsmINLOS4Yhhmv1ecuoxN6dP/wqt693sOUlp3iJqESdr
1oVIT53JtGXHlQ9YzifoZQQC3ixZ/rXPzSMgkoXN8pv01ifsMn+XPD+CxdsaVOUF6+v8omxkAZVc
m88GDthVqx5wS+hOsQsbX7hnN4I6l3HFdrN3LHzT4djf+chkIoK2UTRPDL8xDv0ul3x3mrjnbnl2
r3/qE8qe/9PbuVyItzs77dB+mTgtxdEY1wg3tn6o/jXneCeBKvs2NREAme6Hk4YKn3XTpMkfEynQ
9wgi1Q05WUic1WfoAK31eHcWtsO+GwlIvHFL/HMlOXna4a10tTM4+abXIZYgbdEN2MblF4x6RVko
KZbGYJdycMS/hWhAvKX2yxl/QbLhVPrgjx9/aJkB0wqbcDFKap9E1F2NmIazsPV33Q6rYu46Yxem
RZ4EwGq0aJ1iIOfoMbw67jFFGnaJsVVbsC1cdBc/+9bZZ02uqxTZsCft3CKZCtEvvZsiaYSFh138
h2WKMdcCi+ydVMnb4lzv09gX+toVbQYbO3M5o2yiyny6K3dP3eEaVhP9mV3Bj/S/STDXZR+Cj7TY
9/071CuN/a5vtu1raD+t+zYywIrlaCoi6N/P9PArU8yhNfPSiX0Y71uJ5AQ5xgetg3+Ohdvp79/t
tqrrd34mH8EdHOyYMb6wrwhVidi8d/R4VwNyvDao4GDTceIkv95v/5kSz1NvOMer6UwfnrjgiyaI
ZJ3P0+OyrUm6yBox+fQHFfZprV5iPU5Hl5pK/RAX9I2JtRj9gFMYwUyf0Tql80y1qlHmAQ63B5aE
Jb5m+5wqYDh2sjAJhLHaCqCfAUZUpyKGRo0oopQtml9fR3XUOOGvAmdIlJo6YDEyIm0KTmFETT0Y
mS8HSiwam3Ql9GfIEgCU0Fyzh/TIZjdgpSFRlbfYkTqV+zIomY3m34cb5NqLKvVvPHsvpXMSPgl1
5NwRjvawwFkKrxzsHvVlOPWwQBcELVAuqNwDr18259gWaKY1zBAMj/JDzpSJSVNvmkLRy0OpFh7m
1APXy+RQDne29eRXssaQAZxwdjlUQ0n1l26vXfwM7Gy6wz0kf33fW8NlWpO20fQ2TpxSZjLtfWL+
kZUeUZ0dHwDViuYkb/zhvr1FU/PqKrKVTe10+a7YezDP+LMgROKftXHPSHt5i6reuM5Ssn1qnpgB
Sjkjwr3SWhrQwBDJPViyhVl3Ouqm455zY88dW+dHr3NW/LyyZWw5uGSuEYyMrOaC/wBi+SBGuNqe
yJVgpvEm+iAm2gmqooNPxQDeKkjieL9pyOcO5RnVvBiDOhZNn9cnwA9ei0+OwwGLmtIvXpCDMN64
LDS0BWJt4h//qECHves7EwdcA85VjGR7px2daxNeQVq4Wr7sP5JW928JpXH9lYu97Lw9g7Oe+f7T
omxM2d7uQDTXr0Tw6uLyIMrWtz5rJr8CcDviGXVl/sw9zfppJyEiMETcfg3aEx6HVxlCc28tri9S
vpEgZg62r2mY7pnIK4w/z/A7d70EM1anuowzjKiqiw7YtxFLh0vCPJmCzI4mILQ+M8clQXd4/N5F
ueJgXJkIyRCXrRSODbV3IvMcWqdnK4N1+7lYe5OazJ2PUTz3IPfoE8KR437RTSCc3KWXfHj93QOZ
sh4C03nICtdUpRn+XHlRGj8O48bOlOKnNUaWpdsG05GwUOX2S2z1jNj/+PmaoYQdfWD3qTPzjfxs
5MTZBPoQBm365qKzizBCxMZEroDwJWGqHCS9EMMSdo54HNQl/PJTldwEOsokY0dDqkfYMlj56J0N
qlDq5ghIoCgnjIskOjzJsVnzbadxRYfX5M7280BvnUFAMIOwJwnO6umBrZM3pMzS2qSlpv8JfNtA
+x7gOLmTme056PpBf6pVpiZEaPO9hmXOJWzFkd8XPSPBMB594JA0aQsibvD/BRIknnNlLijrILDu
MqkTfRdcD7IYgsfHDIy7mzOovNyAutT4L7/8+2rImWIy/VFLp1pzot3XQDrcc6Pn0jtyzVrEpa4L
m1o8N9+QcA0hWdzYj/8hMd94ORQLwTFbi7k8Z6/o6O1k/znL7cGt1SE3q52juqNuWOrUcqe0w8nz
3WI+M74K7C32ZebrV1d506j8qI+OXKNjojFqJ9GD/VC3e8Yf/vTSHxSqfeaaz+5Rux1uKF7hnATU
Vf2KRzwYT7zXaLLR1dinHO8kHpunAPRN6DW/gnM3OpwAiLa4hO5tnNYISTrSSvrh0VQv/QEkThTd
nKO31xSEgISYjucAML1/6pBmMDU4KkhAumYBhUu36MyX8vfzezkZKNMcf2Jh8VSMRNJQeiGhqUle
kKMNX54NatvAmDJBQ5KrAZ0gQIsOT7QkmYDgKNQAki85oRkAzNtWHTfJpV2IrEjaCidEHooALMpz
DizoCZ7oUdgsnS+a3zmajxtK5gB1orldBaUKPotPSYbFYp0f1fkLLwSHAVePBa9agN2uiD1iB/Pd
jpVKaiA1RkyyIEK2L8+yhy8DFfi7CedyNWpK3l44uEmr6u59J+hljKJv+fxIMDdET6MH9qPPXSQD
uYlY6qiZutTTH/XKb2yNkmJaxup3kuhQl6hFoIGSIJW1rM3gCBNpa3TMSYceRmXm065bt1fufDFT
+U+bXzhARn80WN4uGVOOexjMMWEjRbDW6JJnlPZ6yanzuG3lZZP5GuctzBI4QNnZYkfUvbWcYf8e
DVRRBNQL9QNihaTrqM5m2swYQNya0v6JicF3ldqLKp181KcBh7aIGbfFbfUkE3sh2lpXjYqj+6LD
QFSghtwUBHk+p79FU78KTtCOGmJ87uhAXi+alI+djO92gyQMtUs7r8R32ZFW9o9jPyfI157r+pcW
RWJ9HJ2qeAk/xl7A/JpEGSOe7AsDWotb7oL3CDwfknbLoJYS+0Fsr+b3PC3aqCTrzrZDuNMGUkRt
O9giXbqKGDNIjdL3Eb0OcowhUo6tGjsFVmopWZQv0e8+WQ2biDjAAKp1doWiVp318OshJqKsKn+x
rjMhAQQxx2iO0QEZnMaf1CegpJrgwJxnK33T/663g4CcZyBdpXn6xt5tDTJ8PNe5E+x1sNIGsX92
C5pVuflRP+QR9fnDMTh+i0L80YhCVsEfZXTN/H8GPRrFGNZPL/taHpDRm/1s33M6ZcHxvyOUlTLu
p2kTo1fi175OhrjxGHShZfJZ92KhN6oX3l/3DZgphE1xo1+MZZ6TqARNZxE4gSDPzOo8uH0wtrd1
FAjeXf3zPTpkXCo1pkFYXUz3BmRb/vf3hqB5rnu+0NJRQAs9DKFc91sRY5cJRlGOD+xrdYhanPo5
y5N0eyJWAioAbOaLxEGws/VOKfLUIWYfgIo1cFPBsB24kZpsGJrommcCcoVtoRB4SP0X5wuuWrjP
q2JG5+4Df3bakV5DK4CCHfxg8vQuSLfAco4NIB5bzw4D/0IjLxuDBFsaqDzWsKdfBn/fUInhoW9K
bRxHGiywFXcP6OF1aWM3Y5lRYL34nvhxkMNc2X6A+T9xBNqwfdj3Yf9ZuNbg8ImNsb78T/iGOVRT
UAuX+8XWH/7Y1hl0Ttnq1nd3b8Q7sUji/OSti1M2N3sHb5pFjKM0SX5gPOJZibJrF3XxDU+OZ3bi
7ZIJXrBE1zitspDq/lrApRQ+PgJYzlWskuB4qtfLXWPVps9m1VnnzsblPssGQAgTP1TiY5zmp2Bo
lCVSep/m5bh6pKwFK5jPuI49vNB33AdZhuZuZjlQsvjWfoQPju6IkeEDyUYSinkCvvq2gFye+S0V
9Zm7QmmTuz9ktWXMsOBPJtezlb3I3hofCjgJCld/ZDapIhIIXGVpJ2ejKvwV23OZVXGwB36nVVFL
BI2t4EA8kfV6jLVtRMtbrI6VHaJy4WeR50byxJz+UPCE6oA/RbBmC4h9RIljePtNbNYZLMxYlTfR
sED0aoRf0kX4RU+pyaVCGSFX2jJWUtdS51O9XQIv8ne/hAbr5syBK5EOZ2l9+/I47+259I5nwNrY
uTtQYGsEF3BqTT/29mUX3aYi/tFapXhkxIqrw+3848w3iV7Fs9ma3AmRS/8NS4ulNX7GiHbY9WM6
2YjYqGUjb754yhUR1NbJQSuuk1Ct1Yez3Qu5RFHTs+bjj2Qr2K7P+/pFKjSAOYWDJHnRInj5EOPN
xk45vGG0RkcVkOio+7kwXr5wGq4L8BqJOWAqnq3zgy5aWS1zFQCAjRq4D6mBpjnGQHdsStxMiGSC
huLXVsW85j0vef3KYQDaaj50HJJB5GoQA7cAEjp+znB0klwIH3SRluwSA7f15gEmbUE3+/rINnvC
2LSjHGPUkpK0Tp7CtMv191mqSUXJjFpLlCs6MHNF9ySdHqngd+duQGdZebo54jDFj/71FVMsbKWY
8HIGqmCl3xliK6HuaK1mbh8mmwEddoXsX5atwJ24wiQHJc7IYm8AhHHuWGsaxfEOQ2Bl2TB5DMZ5
TKCr7PQSNw0qqMMMptWPCC3IUS42v+3pa9uGajwUG5ETRPamZxOBqbpkRLMtEZ1IoNWeVhOGmY5G
pObBRtqIN1Qct1wPiAeGMZ19gs5qpI9zGI8cetFcaIf+DLO7NBtMkx+9T0W6jpwROKOkgCXG8is/
IbNH2O4xi2ol178hPk5wXGnjvXNRWLbXe1fa2u6xKttq3bs/QW/fdMEt07kd5KY+87Z6rDPyZE3H
Eq6mhY+9IHtIJxd1oYZ+y8/Cr8nFqnl0v4X1mC8yJ/I9HBHPY995qgYLOohwCfH3sVrlOCtjnV4c
2H6zeydjxrMnicYKJcdSAPp1jK2FLuSX28VBXFYsNftboooy75T44tE4Zx1+guL/3S1tUz5L+bvY
hS61JiCnqDHIEeKt6Ep3d1HNQOOfIjc0jF7JDQU7QbWfOsa/l8pzcKiSkCk2UJIk30nRyfJ9p6WW
Agph24+7Y7jaj5weQOp4h7aeSeuOgv9T00pb6kmCbceV+9tPQ4yyW0AjHuLAbQYOhERcrzthJGzh
jWBcLLGCRhC1ZWS0WQnVQ5H40N39d+sxgwXTRY3LqGwEdlNFaUwli6URN/4TGK9/IfpYmd1v0J7o
X5RDo3f7UZDyvNL+J4pfDvt1SBuKIyzx7jyeqOuhbkXyirkw3yJCDQEBC/6RKz5zBSdvbUXjFJsB
G9Ujst1xnO+H4JRzbFJGJ0OP7PSPll4I4X1/zJx//z6cx0TOT8li9c+dAAq816ApIA8R/aJRPq7I
rP/ERr34SYdtF0cf/gtNcpzSzlV+HfyUcS46Kzrfm7f2B/x8Dp9NJ0Qkd/gO/Z9shWc8A8bXkxsC
1eGQFKNNw3H9sB/exw57MOBObm0QAkYD/xnrHCco0bblGn3O1pCUiEwstGIG8wb0m5ZPhGD40+u0
FWSCOiDc1BShPm6NmKzosFhjTDaXB2PQZCu1/bAfeha6EldhUkyYcncCEz29g7fPDn559yRVmYKb
Q8071skrLx9mSivhExlYVUsbIOC3jabGiCY8odT0oPKTTupGB8MCVKoHAid1RosZqYCPmjpxvnVF
bqnuKV1A++Mbw+1ddER8o61jG3Ju4xu9XT4i7xV7JiffquCpwveaQ+VVzAMk0yqopT28IGbl6yvY
L2aKDSRJBltVtmio5pgkSafxMnBe6GJ37RTzNwgWEmnp5L5W8VIScnbFBUX0OzY55KijYLsia7o9
H9H4fwJJuVV/1vLMP2aTHSi0URuerN+37CPlTtoPfFyyEkCrmjLN0oiKL0WFmoSun3h87uCDQ07v
Ao3ZkUGCobq63G3TV85mwxJfxEosdcLNJjGUD+yD0PzX5eHm3nEpJ5pmw872MssOzDizU3UBMzPU
nidj5xwMg9V0J6v4JyRnxLg1Qcop5rNBmwTQGwkWgSFVkHGb5CuSvq0by/bYWpBGWwf5Og4bXYoI
bGu55IfON3+Bb5uVIDalnJ5wLoSUk+Ayk38VTr/Mf2QAPts1/H1K6GVfRKKFFYbwW8Ig4EE0+8WF
epzjhBz9zqe8Pj9erduNVbw9tu9bypDBQN8M4+nTlF+78eB9u9Y4teBux6E4cHoQ3XXAvjUxv07+
HeaGtHkgcvi57c6U+HmZmrtorvOpt+nTagSzuNn99d4BFzFfFWB/9ttqaJl7G/BYkEWICHxeqX6Z
RPaYIkG3E4FoAaNfXplxbV/sHkGiYMim9wJ4+FagHkJJ+SQxLGYYO37vQtAQ+PmPDypX4Fb6czeN
IHCoZN0J+YQW/UF9V6x1xk0lGUrP7gqv66/wks5Br1XJSVLigKAoUuE2DAD/22+otSE0m22KKkiW
NfeCVzJiTbO3Zjkhn8pGUD8nT8jCXLxYeb04Hj161ePZeh1DAO/ZP55+MdY3c50YzETkZx2GzXW3
EIpNbZEKGtQ9LAHE88wcvNW7r14Tm63sUltcgZBAWlW948BUvygE9K4mquY2/CvGbX4Ia2Vi7Pv5
gXVzffAGvCMAL+GlNED65EbEMVmm8t1OAlyGcJF6+lKsCJBmYVxr4PA2b1vf2ppGoRMyNHqMJPTE
ORKdipF7V1pqIoQCG3FuAtgev9+8+HnnX+tgrmh2YmCr3xTVKsl3i2UWCH9iPzsb2ughvdJRVXfS
PcRjvERXMZORKUKdBwapWEfhDjmVIs47MxV8Q++xk1SKeJBjTZAdEnCXbdm4crOoVHnl1zVBmUJp
0QzaWg6121S5vc5/wU8uyrM2Fl9iWqyQvMT4oQD5uu7dA8apPnVmg2oeLx6bq7pfDjZaLZHouYzk
2KOra3D8nknIk8qBW+i3EL8ACmsqnoqhFXsrXnig2//q7di9BIkC8XF+Z7tyqZOWJKdpznTtJhyo
0sI6oytJGCPhpceA+WqmSJEYoLdaOhnx/l/hjIWFJm5ca1rbYk9gMnw6a9SVPUJFzl1RZjpO2DzY
+KWe0PW2RIN2++Z0gVueo9oDPy+HCH4aYLUssS/nn/IPycjuyFGhUXE6eDLyWlbQf5yEqKZqM8Qj
RuGhX2U0KlYBbb3oRqxICCCENOGqV5Gj79JGckWZfDbTbQQxxP0mEnLpBaVlVWA8RvvH6iM1iSrS
2J1js+f0tsKm53S8pdh1n/7aZcbLs4LUsMewJ6SZgsoSOmlcQwbuQiR+tB4aRBX+fql8Nte3BN9m
aTqX2DSnGgnay8TWY/h+UfhhhYvOviS3dZ3FKJWrkusFe7hXqm3Dv3QSYo86Ey/Otpg73dYOMdS7
clm5914zrMRipZqn5UR1tf42aDbRkw1WXBDOldvKj/m8bJxBNFSBtiRFD9FXjGRLaRB2oL0odMwD
mGPH4Pzs75oZ4LSeph99vMhtWqx3kELVWflVfhJlXtWY3QfJnBp6VrhYkvuCEHyypSNJwYEqvQd4
ZSP13fghH0ZLWfQJh0OK/E9hyV4qSVMxGj7vdASvNLfcqA5ZwD6F3COAK+jZVVffZDt6JXtcOD8t
zmvXbigxjMqEXOLM7jPC5c29fI4Ni8Y3bS72wnJLxncuTJUzs/qnuMn3Rg5H06H27kaXpRiYICFv
XZaWIsu2rso9C+6dp1SUjc6/Rj7sMH/4DkfYGhMvAtUfnSf5miw0JKcjvxLOEzrYIshqdHYWSpoE
tWf4OGUenxYNv5LE7rHTWYDatsifRif/rcqi24lyengP0RFy53clIlmtlL1l+b0jdb1ZRxtIQZIX
Yq9sbw7DbU8ntG+JZd/d2Dj8MUgCE8ffAzfnXTDYDxIhVpO/SR3t/SHREU8HybKsK753PrQ/OFOM
zU4srzT6WcTvNra84KxlXNpf5qmV4wzmX+GeGdpTOMnqGyCdZBDTEpZK3fUnEsvnCZjf+yLhx4/p
B8+Cy0qlLgEzq4/K69pGWnPusbZHyZzTcN4LiVD9gSIB7yIYFJG4Kiey22nQF/sMnBQ8IxMAlmUp
uiAl/7NTXOknuuZKFq4+pzVfmAMGLnVS4XiwbXU+otaHL/1TLpEzONFaW8PtQdeUJcY1uWjsnsQV
awSuqOgoTXQDbIgtXwJ0e9i65BlVO+ONGHRCeTwAU3eujJcm5zJdOH+c4GlHkO1jEwby+F80286d
pR+JM06Q6xY5d8wnKqBG7XT5G03OLjqqBMkdQovxHJww/T5eZ8jqIzy8wCHQIc6knRB6upvGitMM
SbASvwGq/BT/g2rB46GCTwFN5pu6HeMfvGa0xUotQ143ACwCuw2+MNQxNBIuJgES4qKOheyWKbU2
nqfgsJfMCaZDzXBlQIHe/D8LLaNFV8nIfeijIJOnGYaCZOT8fkKqVI+9hhktTUk6TlRf/cr9seF+
PKcJqZgSg7tkHafogxmRLjYq4ROG4ZPfsPlCEuSweyIrOhEJ7VPNBbVd4ig6x+rusdGeLzrpPgKp
NgHqZwMaznYyuqqFEcxhkoRS2JopjFC3WoQXTPoA9XSmriT7odIc+JeHkQihNkp/ajuIYi7/gcHE
8US3jlMPhVksB/j/tu6mMK9FCDttnAslbT9obpXUbQ7n7eUyule78R9XJaY35uLvUGGj/HS757S0
SN0GHHThfVMwf/RRYKKXGwd3KmFd7W3OjL5NQlFzNtckXQszbbIYXIJhwGwLOk8TquJf9p7+3GJs
7QXGy8SY7dwCGCW51qC2Hudhp1PlS5KFir9u7nJQ0CJuBabj5W9e1lrgHYXMMig9YaBmd+6Z+z3+
H48FN36EGw5v0tgtYvLnMubCCytQN77giI7sy4wyeaoz7n3vrDdFt22ardPP3InyMC4jaXGFMm0m
We2GZAOByBX0kSrJxfIFm/tdI74CPYF50lGDON1mMbAniAZBSE8cNjRJVGEnpJnnpzDnZlXLkD+/
ypQ/I0qkrFQPTsK3T1ttuOaZPm9IO7s7V9VCBOomKBMDGaxsL+VwnDa95Qy6YvugSRf752snLjc0
9X99A1VOjHfF9tau/WFNKTWhV+VNQX8xmQ5wDTHTs7G4FqiOnDOWnK3hGr5b3WLT7TxgJIo1ufbM
o74t5M/OEcRLFaqFj+GC9MKfbTxLGuP21amDzcSKX33hQHxow6eqLifdwsZQ0ZpfvNCYIHKsLQyZ
2zn6AI8YBwR/vy9BgA2A66fyh2Up6EXWf7yjxwZu+7vxL7iK5pr6AAlPWe4WedvG+Z5+2WExO0K/
ILnE/Y6wNFmgpskxqdfHC0ssMUkKJBebhVRjIdJNUlgh0H9at7HubZs3Rik4wq9bvczT0ppid5CI
8KmYZWR5lxoFoX2qpbVFhlFy9sBKNUs+4ZPzPCsAEODrcpx4dQDLwKkyYrKFveFee5gje91y9MTp
fgVAVLeveTqN5aQ5azTIr+7V6tkbZe+KvbJB+IzptvVJfhbaxlIoKVAEvPxGWOv4haG2ANg8Whvh
C2gzb7feTKP2L9cY3OQBQjbSUUWicUCx0YMyEPrKcUSw8CVPBeS0NyNigyWS/BHu2HFMdu+n8S5G
/eqntQ0tKpso9Z6sjz1XjngXrJCZmrXKsGjY5u5vKv9Y3ITcryvW9UgCO2PHN9jpNZ4OaJSKGbcH
df4AXlgyUGBFOOyBloyI2+icBdo9VBbP8iOETe+fk/c4WUnnzyER9pgUmW25lbHUyy7AqTtm5awQ
czjcDE7x0Lje/5BQfCtaxNychXiTPozkqkOxvgtdyeKC1FkDR6uRqUYbaj2LlBcM17xzj8y8aLD8
lLqgyckbAC3N681JY3gB2LF/ioWWoE/BpJ+VOseqxqeUkrpSTeV79cOixRYZhZG1eoKAs8W5Il8Q
HqPBDIXtmGygyXzRswwHGHyvF9fiIdOv4oUOSJ4GKQ0qEfoBQicBu1CIy4Oi7KWCrRNCrZFGp07u
4IsBoa4iMuNtoWkKizQAFDUQXjBQQcZAhGdVwcKXpCudKYSajLYfDB7qFSQfApg3giBly2L7FY+P
YKZq7ovFFikhKvxkNtcLunOrcs2BMAy5NEuym811RjYhN5Z+2jyUItnxmh1QWYldm2AZ3qbp8nbA
wo67WGIIYrVYOw/Jyy+7uz9AdqV/y+PoWKzfvamEUm7cY2aQ+GIq8aRJO71+dSLe7qzi3Eas2Lhu
wZmGUbM/0JJj5Q0d0g8AKpBO1hBRUjANqsXUei64dbYLvGWzfgbCfZopvb1PcLVbc84zsXaXhIRE
bqTTC6fqPyL8qwL01Ia1Zx1tLrfHigRFfvaiataIKjnrNn6oRmsouGRg/YQtrXiGktq6CaskBGZG
U39Tcd/69qWtUmNzUVpqafFCqdMRvWIjWsGB3WoHdmb3bRuyCKE4Kmnv4mQ5zmrYoc4QCxI8NG+c
xrklnKAEECBsqZWAxabnutxeGxDqpXV+by/k/J6oj6qtyF+tHRi9kQt7zgt5EdolPCV2LTLqVFN/
PQwXJRzZhp+Za8NijdHjBIB0yGlQ8fnVqGvchziq95t4Car9My5X83ca5R8XYcHSF0AEJZ9eS+hg
aWuQGQzm30UO1uokygLA459hnd4mqjeoBkEfd3sQb+SfgXGwY5sSu+9D3i31MfUWVU5dv1sL9XKC
NUaPDFBnyyy5hNU0wWX9KyiNLVpKr/gbayi18Q9+250uhSnr6qTcMn4MjRhJs2RtxshdePCV9R2m
Q6VPe3ydyc+utBaG7z31vQp1K80SQXT5SDEgtsQbHCvP9SJ/2R2R1f24w3sIsnpvt1tG2WUi/bCW
1iuojfAYWfhApmPr/NdtPZZsupEMnCWJFgXYfTbHcIiNhij69pNK7m3Dt1yB08sB1r2IXI178HjW
GfFkcIXKFOCKEMn5T6xW/Ywu0qMB3+xHI2y5hWO6xLNznal4JBY+3M9HajC053ej/sEnBpP66tUM
lG88BdpjLLty5BZq3diZ27E9k3olp4lvJerlBO/LYZvDJzfpzho00tVnJxX2sl35vEnG8Tg1fIZu
YlenlfN3hquQqFziYaFZdpIjx+dva4MCzemECWIui7FJ/MT/vfFuIu+EMHlVps+doJLwWPttI1AJ
Jx+Gv732+/Wi6GBG3NlHeuRvA3ZCLt0QLUt7H3S5uL236dZqDoO2dr/v9W5ALe3a0ltW//Up3vBr
s/vRf73V29N4LFqynCIEpfKLxMDPg0ftdQMg5bdhBmSIpVZyeamhqITV2DZ0ZtszmLrWhmfQ4kv0
SMayW1KjNJt4EekKK68oH9v19u2gr+PfWT22aqHE8G9Nh5dTMinUtwb++CCuRHP94ybSnyZ9e1Q9
0CMFrR742QPXOqyTtrI8hzvqefYRVvjBcd3vdYjPZh5/8bit7bxBeYK9GGpLyYTw0RQHqP9ZIO32
gZaSTixiChxLz7XvoN6dZ2/kwNl78uYSflSZMjhC0RYO6rQQO4AM1LRlbFsfrPSX+Igt6HIS1+rt
kg5VmxcxOcfBq7j/6FGmGfQM9kz17/gO9/knvd8lSV0C6mdc63e2/QPQGeDhebevQy4ke6qiOOu/
SQMIolxRq9mlD26CNW1G8IQ4NqreqoKwuap22K+AdXxSWr6tQ/fCtqjGGn/Z4gpLndxkxRYBnH/L
3Ehi0O0PyiMkm8oGr0s3wzx8H4O1YY4gz2JJTerp5bx8IzRkw8z96mENr2EII1MMypWx3XiefvhQ
04qi0MOQpx2RyeOOozNKcWDdhsUW0zj8/GzWbh6Jq+2D04I6FQcAt6JhgOhucER3mopmwnmm8l8M
GrNb33esnxbJyHyaZFKn7ssGvYancL4qDyU+LdufeisLTs5x8yh3P/sEYgHa3skZJbU40s8LNNkr
gpn5xKoWLI7pV9IxbH/cIRbd4G/ny/Cs6XnEcBej2RErB26dc5DwsZDzXBp32X1bbNqVwy9w+jW6
kNMD4xmhkHs+CpepFrm5QcqIvTW1f1A1azzMZh4XF/x+TL3xStqrirHvHfp9Bo8VMXfHDeow7SB7
0pwOUY2hKa0r+ToMqvxtym9qvAkuPsT48zMvOAAfVnfejTNDfDNCKyThazN7685MoPyJG+V2anp1
clxRQgw5UFaJUWUuK5wX80yg4V82VMNH9r+q/F3/Q/lPjX6JV5UU8j/I28wXhna02adg80btYw7t
mCpHOtfyh/qzVR2RktL/J/DwUAb5NjR8km81Pp7zEtEzjeKCzs6dduftwc1/LUYjIi/1+mI+sBSk
nCkWD80exa2+hwXtunh6sDOpR9CJeELpiwxYkjDL1QLMh65K9/CswNFiGhJxF9nrfjuy//8MIaIu
jgs8Gip82Obx5cxEgNxHda+otpi0fOJajrf8fz50l8akepAndTV4P5RElll/buJhvHwTxhcwYd2m
WZjowiQvTBDsSPFZlSpQfUGA3qksrZdMKzf2cYCB6r+XoRMxrkRRy4UPlyIftuILGskAPP9uYPuj
AQWctDPTtbx/JtmpfJ4yx0TVTa0WZ+8q5OAsIQHiIUT2sZ1Adp6HGaWRikjKPKOV+oj5WiNHjVdQ
Adgud3QFe0O8RsTb02O8+dvhsiz+waOnIMyS3WnwFUCKHqUSrRgDEeMTaI+fxxx0kzRjcGwRAmCQ
61TETIlg0bzjA/xykY3MpaPWSEjDAlVm++35rclKsDiZfx+TVgO0ZiMLRc7vEn5spLfjK6TcyQHO
N/bXgBR2WJT6PxO8uXwuGukQvG0XBXhdsV2P1ICMSr3MCOAtDNzecK+jHv1dqcKUw1aL/SDpKlhf
UoKnWwwOsO9Xxtyx4MfMDKgk2woH4s7bZj3J6gDFwIHUfzXw/wgHuPKmlibwxd5G1rp8VRcp+YJ2
cofAfeHHBhvmMBMt/b5M05wR7dQE9VNBpUs3MAwfl9CBVlQN/Ub8UJJJSllAjnRqhCBgTVsdo/eN
FGa79TBjiNwK6Ieq6zCqv1DyVxjw2CgLr2fvXrRdfTbb5+U/EV4hPwGuSLBzQZjwBF74Mq9IU4fE
6YGoOpgMstRP0pXnQpkU+Oaa0uVxARvO69ePVxAMmbnEtG5JYJaDyafoglC+EHaQLVz7JdXMugL4
lAUa0ilRiiPeWjYQ0fZujJHu/biWHWTXel4E54fGVSAMipC/6DWoiVbAk7ynk2Kz8wVsX4aCXNuu
g+bzGwD9GNka3pEQhvt6i3EseY+rxNTeo/fW3gNhpBpku1sCZZQLik5WpaDiLLO/U3B8nZZJhqp2
8CwYt6Q72RVq6g7A0s+KWu8dtQefZl8/+SmR6csWxZlwZtkrq/+Ovol9r1MXFHswysxzeWH65aV1
uBISloAtMmGqI5v0B+OMgEdAjSeAInLMUnnZR0dyMBYLdnoHJYmjbT0l9Slt2AgR4a/dEN9TC/MG
bNLp7hfL89Bav4irfPYI8HlGFDn2TNYhvT8qoqjbzKnCOy6Dnix5UZl+NjQdXZxuuWsP/vzHWT4D
HYz3Q0YYj8liSbYJwHsoiG3E9UQgl2TyN7k8/Y7j61jOOobpsLvtTfRWEg8sD5g/ZEugwqeI/XBI
fvbyGxgrbQFkpdAupu3H/6YlLWOjNdbUY0g2I9pym6isYxfA/q1YInKpfZRRSfoyCS7rUPmExxBK
p4aTYdaW/MumJ5dmrG9rkcloMWdq4Hhpl1/L1D4+L0yu8UDGXWBpfPeDLPDsm5lwvxvTBCuZYSfy
TCvkfq++czevRrXPnP+Gft1iyb9pSFoPT4jvnwWRpgVJU/S5qk9M7ZUUHQL9SOZHnepR1vdaNYzK
ckFmghS4fEjdqwK8PVZcAEXH3lJo2dqBCyRXMile62/oKBjYbuDgufHauCKViktsXSvDpvaPySro
GOlV99BkqubPHS2Hz7HZ+yAl2/Ool2k0LHSKjf9QAfsuXOqexR/C17oUqfzXxVfswpcO3F+cIax8
XJH+6Rour0vP5jiyJzp1zmoEkybJKT8iG++rZv1kscsjX6euCvOTfHRDV2XhpxdWg/VR5wEfsxPP
6Y/W3ZfASJYjhFqIzPbLgbRN+DcYEzcuwpxm7gTSdHUQcCzefKD3h5c0bjqURuj+ut4xbXS3mGAi
jJBjGJZ/pE06Kh6Zq0aRSOzWFCrCqUzfza5gVVUehWNx03tIuApBUVD4YcXCnIfeoRqvAMF4AGgV
vp0goBY7yQXU5ex1CKAVbkNPwEIa/BgVOogQoCbPGFXTSFllEgubF2V31yTwwZi5l9p8X96h+d/n
z0iWFKGmasJ6LAPD6RtlPLWVbyzptOTC81EUvrzjkOQ3KCPGCyFoX2uWoz793/MZMjwsoXyJ6JSD
sHu7uURMocRnCRxqEA6skF+Q/yMRwVuAjjcaxFljiMZ9auehjflhscxzPsLWHE9Cn9FtAROmt1Xe
61igstngXQu5itvtR+StKPfF83EYe4A9pB05bxsjQj0ddabjDz8tJ8Wp2hvg5ptBCsgZPTf3Ob7A
/NXeiStwx0Ps1FRRwItLj8ORtx9graC9QdafPuVA1JjvnJn4Fb6TQvSKAwQoe0Df9EbgVprdkbIJ
sS9Y8WX+wncvJ+vQs0gAmr5ckHRLZsTvjWNry+oqsIGqOQIX9GNxUM+YPw8RwjGvsqHxXIYICFXo
ttu/rUTnJQJ9uAPKsK/85VM9lpw8dXWZHuFuRlfX5lNy3W1XIV/iwz1A6uC2MJOKnW/6NKFsgrax
Vo+xI9WxbwIemc5lsg1cAPovCdskgbPqXkt8GjvphMEmRAkCTkyG+7cXCmJ4BBWIM65zrAUPXMPO
tBkQGs1FQIq1ihMg9dGaE68ZubhEUFoa/PCQpAI15ZX7wngbT3DlMhTeOK+NVc3r+IggCrMr4WfS
3rBVIBjlU0Ho3bmoRrQN/9A72n22xTqL8r9DYUM1ZL2GJeibvERQSiTKUuqvl+CLli76ZT89+nTp
Lh2IJJ4j3KFWTXcZXC+nRnxcd8P41jrcVFNgIfXWGn/p07CyBh25HkQqXuPgjf7rEMx+24VLoQ8A
xltYVJ34widF9NpwXrRZRSDFefzzXuuuOfkp3QDGAjKgxkueIExbqXY8vqG+bqMYtm6kZpkcFKnr
SdbCAJpfnoRGla1G2dRTjNyWqODUJp/aODELOLRCy64hVkadQgFp97jJ5NDU57g+jS81GGvCL+nh
8SeGWl5GsGB6vGSAclzJ3Ng0r5S51HnXofJIRjY0ZvEZ8AfZ/NIYjLQtQX6Ne4g9XAEvZBGft5vN
E3bu2u4wf39PoYktlnvv/3WYh1MEdooLqFawe83FSQqjgDyd9/SlkOD6pn9gqRibgyjQIECfd43s
B8AOia0Y4rNc6l/sqFGda27+CG268uQZq/CThOjxF7q4Syq8heSGTUgcbU7/GaOywAVyx8n5C84/
5yBtKjX05Cp8f+3oDfCVS8+DOwMfbE/A75kVN5up6ZpEgI87b85FkQciFOpC8RkB6s3F9v8ySvKo
sj44PeYOq+9awiXRe4m7ZxKKJi8jgwNGvL1UlVtbFzT1oemEoRnvNIJeHwy76Gb+qtqFO5qeJQcy
YwTZB0peQsoTQipEKNav7o15NOIR3MDj/u2kIJ/0+TjsFol75WPh9nSNrWbLLGLrY4SlemVihF0c
8HTF3KKnHBEabJf8uycAkDWSSL7iavmmXtQnl4+xUZVNzVrDxYpy50y4f+PLTy97NQPhcSDRBZQG
lB/IR9SA+HW/qVFYKv8xrnwMKga1fAg8Ld8Jb67g5L7+nKg/8A25/0nWmdWH9cJXue0/gWvyXWtZ
YcFVj4cpmC6gBzFAVoPtpOepmOAd6wJ3eVdpZ+WHy7ecqYKk7NaT7tpYkJY4/f73JEOADDBwDVco
PpkVRKWkZ9k7AvUAH6vWt/kNPf9liT6UDI89rQ53cGEOihdOI3OVK/ReQdZ7EMb7ot+4IzqUT00Q
8WTSlkU7BOCGJfYZKiyzjeUjRWMFY87WM4zDoSRFr8/9GzENJcodlyGidwFc1kCCU/s3i7Tffwmq
Hr6bRKbIEWIWf2N1MQJkxuiPp5DcQjFMUAL/i5Y4YZouJPkCNeydXvpnUdBojUpEXgKe44U8iguW
7YEYQQp40rBqs/YC+PHxBAcyamCUNl//YTxeNlYmOND5Tr4hel5WglQaADArCzHqOXHub0FupYIq
ERj42a8T2xydENM2Rr10d3bAKiqx/iIYXqqXdxArRVnh/eOoqi2VjgTb/OQtojLmXvUkmlNXH0GV
u5uFEIG4e32HR046HL8dwwGT59FZjY2kGLLl2QJmMGhsez9PCcOe8UKXbh4U9NqPApAUnx9ulab4
BEycTbtljV7CEkK4Z6PBzxwLUFAcAqHgaTUeFi3h/90d2B0OKhajnTRA1V2x1zOIs+/6+viRl1aI
qzv7o2mDQxl42nTGd1UBiYo9cfLlGYQgcWuZhsW2akyS/U1IPU6IigD17BV+JN2SeDvkeCmpV3hz
8yTwtpWrfJwWiEQMmqB3hblWLj9LlIKR2GZMVQ6sr5I+CxJFNITz9a0gDhHABhlK6hoPi1ALy/YD
seEQWUcLvv2iFhM4horYrU9gPaUBz87UWCRu7Np99yZcRuLDL2StdY1+Opfo5AdNm2VfLfik/vDa
CQ0CmEa8gCRdtpfqlqOvvHKRcCR/WNgLPpXBwcUwV+SbJSxPuaDSrH+DEFOPXioVX5PxSzPhLqLr
5xhd6dbqV/hD8HBStBUefUWVcX7cWlo8V477NkNkkgFWCoMpa1dDHrk2T6uUTHu63nLofp8J1b7A
OsK9g9cTpYpaz0I2RpbIyzgyjf3tqU0b1RQrrbnZ15741jS681iJhMRu1WeyRfBVAhgO7dwU55sU
5q56Qndq/2vtGcLeCRVdAbLH+LR9ABhGELnF93YnrRVjNFVBBVe6XQVwI3GDrGGK+0gcsAoNz2v+
dMxyty0Y+Ai5fD3eO2fH5v9fAhi9o+xVfdlN2ZLIBQPlpot2QHKuNaTVa0FM68efZf80nJ0fOMyd
tPbWEoO8UK0Zinrcly3jto+St7DMBYSYjDXGPxlacIzX1vCUHPjTaHXo4n5a21VI1ZXmmM/+8iUK
9fi4iU5Qpz95YnYTj4qfjPA5Bs+6XPi/2z0+ANT25Bfavs+oMBSFyk/U7TKYgWN9mXCvamaOdPxo
KPJE1HId/jXy1fZh4lq/S7uTN2uFWsMP+nIlSSVI3+ecy2+vqb1elt+ig4+KeP58vsUNOAiWHii7
GI8DxYH4kn0bsh/7gJG0iPsbqIYo2XUZPryiXOzUIGwUT82SZ57TS7ERx4I1GngwcghLEQvCJdae
rFLXVMXoiP9aBer5oOpOAYOvPNXjdzpFNb5nS0Ns0qKQ2b2u86+EMZBNw6de+N45K2e4VgceG8A5
2ROrkHpuY+MVnYF5eZqbI2e0kc28XdHpDfQmM4Enf3Vbr0JqvbkMVF9LvBSDo+lhvgrsXExhf8Kz
yeKGBgZNUUPHu0EQQNzJdjSZGIAc0ymdbw+ILgxo6Gkv4BO5+wZ34NdV5cim7UKp/HHMoAzhrqOO
LJMptMyGcYtwiyNjBM+XxYQxDqKvrvHj4jdo3THJ7fUXSCHVgDwzDchrLD/qnQB0fyvxf8zP4YpY
SIbD1+bjrEjoo63dY+WxsSwzLl8eXkdysOl6EDzYGgIBZzfciKNvbir4TS+oagkXpYTMxwKKyF9H
frPRBv/Ci8gDU85FHYD2/FRNf94yWZrTSF135FrhLv2LMEo0c+WzvuM8PxC8nbqjaTVsT01deu01
uT9/QKURhFVtg5SxN0kNOIBNwCqDb0rOvku+5xivvYQq+cyKUa05bZIkMwE++CZcUPVbxpL11KTS
groImRiU+SHPF0224V+bTuiAyzzQvzMvE/f4A2WZ+FcGAui09XD3OpcjYKBBq1GxEcVWLDMRXnc3
RhVB/BnCMye1EyAAUDUQftiLAUU3Br4H2OKBYwXGADJB/nUUMXIMedvCuowr+bjtJsDLPsfMRqau
f7QK6RC4NB5TaFRcT3QFEYTd6q60H1osFHibvmwrLqW7bp/OusUhZ4zU/3+nsQ0xb/6unlpq3sG6
go/hJrS1BRlQUJucjFrG2LzMEgER9thdtiGd50gFOunVu6qdjvhRDqptKfy2gxsX3ANFNJuYd4bT
dls17GqSKSR/fpRXWGziR1UBzeG5eDTYCKRImk3UZ7zgUtZnLF/s8ypd8T/bjk7UpUsR5PM6kx8V
o12kkEiKSRZHfNB/JSt2xAq49er23Qn95fWILWQDwyLykimKAp5kOCZCHZ7qQAzat/Qi5uwkexl7
rszYY4bqB2rrRZnUctSmuDS4XacXxVBPdshZtt2PHzt11wrfKfFVKNR8PMFe3QertbfSgvKoridQ
TIk8IYpihUkxJ5WriyreOoXcXEhFP7TTNaKGCx++qX7c/cr21qFTgKQVRYdEgKkmueZ/s4tfyV/H
wSDhNiCFU/2EftAvuiqTZoCpeYTypMRCAkbzZNJbG39bvyubzmINQEp2jn/a1lUgefFod1pubfZo
FE8LTvYFH2thQj8JhxkegcpMBAbfJcUiHF+OMWm6EEaa2p0YL5cATyvyQ2YGXJgW0GHLudjrTu3i
LmIncRc1BYqWkGbLAF+r019+ZXyOvCNvgFl0a8m1Ll2CzZh4U1wEvUinM1BmkK9LgVf/RXZJWXqD
1nnQlzLay5BqCToOJTx3QnOsejbEK5PLVi72XQqmEdQAuhDTHxhuloxEhqEpPahYCNHxHGkFdc7g
RMLyQasSfMh5XKdlPuyrA/bK20cTeoktTgI8dzCSZN+RxvziyAc+HTfv3qkGhm1F8X2sD5zDq96d
plutMWWad7qVcHDV8ZWZNCmbauVzDNsk4h/F+YnQPtkOyBzmnV1zDxJmTidjzpVOBCbSI4ouft2S
1Fh5K8WRSX/e+gfdij6wX6SxBieM2NX7nPCdxaWkgxETXFh9dFLiblR4ROtNp3XDTgpCNzHaDVcF
3K5XS5sjEEG6HEloQqlUPLXVCIQr1FXBnGDQw93FqK23cN4dsljsdhkpp4G+muoCdkEXlTqx2T6Q
51LxQbqa4Tz3QMblYh/PuaMEQCaFfZRRj6OhQl8+7HH+m1TjcH27FEMpg8NshlmLByKDAXQDWKBl
y2q8JcF0Aher58K9/SCm4mdGxueh9gwvAzGX/an/CTb0o6WryBV6O4zBp/sKIJ9oMIF+BXaBMt3j
xV2rgd9EW8lzh/6qOgF64OF85MHXn7vgAy9ZUZqeJXiCswJc6BXqYkJFDq2QRr4Nn5AG+4Z8Q5eo
UCMAKhLwd1QaOIyxIbq1BrUufCIl2Q+PUX50LpUlXAYfeKOrlsHgsu8yRzsIsazXXiN/roB966f2
5/uNvkw8mZJrsE/h5c3TdbQhK4sDpaYTn6p/mZ5ARNwe9npf6eVHakiNf8kvdIGwvT9MZBffckWK
85zWXHusU3Z/ocKkfQ7x2KCooIe7VZL0ayvEfz5yYz0dnQRYNBmm4ODJA7dWDp1aoC+Zd1wAyBgn
711zFCCRbK+i7Dm72IOVHijYSe4WT2I5qTCSl38bzR4plgl9AoJ90oAzmPrOUUnfN/8Jmz0troMA
Fz1jQqIf4qlzKf1tvRfWT00BFwYZ8Z+ntQzPOQ9sk05vRcVbIxKodXpl0QMIkNF/7w0aRehWAuuc
fVqYLdCh6sjmlZR/jOe6avdsC7IJ+uFVbcIkGvxRykwnGI0xGMfiFSLkes5WeSQ2HUbfhndQB2yn
S9rupHeeTtTqTfF6Z6bnfekX3tQm+Ji2mrsATHGROU1RQmvPE5L19JKtLhA+p8DTj/JGGyYZTpnr
m9lYx2Oqa5tVtZD6FPsimi9LRn7rB2JDlmDCuT2B2Tx2Mk9v9LnBvESc/WA0hkmYvI+vj6OIJsPs
YG0eKtA3QU/Wl3htOkNbqxledOESXAjbIJbtDQy6JI8tUQLKxsK8bCHG3jiuobaVe/mKle8Oaweq
fSSG+lZ9IIvIKOAIHE5X2e/uEoZiLgeM7RomUSllPQ8+iyXdvMqusZ2Entcw0S96yBlgjSsm2c2P
IBvWqyh7pNZo8knTATCRAg21Mfd/xiInBdPEOFFfyNfTNf4wKl+4dEoVrRUuAp6jFHIHrdCCkMBp
X6WhZJjnQrgZsqIIuag34xKk3+oFzpOHaZpUhQwPkc6/FyaTjMsr4venD0p4wTgV47lVhIajs9R9
5NuNk7UVs6OhwPsxKG12gGhweW6K+3hQmKBh4+S+RKSTpz7yV0rbfgy6LGwE8h2rIVl20lm+fN+o
ZJf4G9klEvLqQ0rU33sG8hGWY4nvKIOFjAF00X6xqpfs35BXOfrCDQ3oOwpVnp2jJexbhAiqKOH0
a+SNUyWRlZuYUISQQ/lOHiWreJSib0j8+fUnBl4QmVVrI8Ceo0GfLUXhBi9dhvC1wSrn4igh6ppV
Gi+WJXUTB6rHCPiAjEFDhDKr4P+sGXqgrCz7oRQvubLgpqFzVaMhvX8bCs+kp/9NQ04P3yjuqdjY
KQt8gnWlkRIfhfaE3ZNGFOxPbejLg8FpNFkqnkWLFCaQ4ek5rsKRZx5cSrIXjQFRD2DjD4qq5MSH
s/756SY6X7Fe2wGvy0Y1+epgaRiVEsTgtmSClraFATfZ8pE99hjPDs1K7HaRBj7lY3/hDKpvs+2d
RKRQ7ueYcQwhVeICF00jcsbeCYHWwk2I0NywL6x/FkThqm+Y/H7YTEezOxwro0KV3b+F8KnjP+cM
90+HpdsnVZl3UNeZk6SXRn18ddOvSBy58Bdg7KVWOWWvXKxi1OUBzwTnQPU0O4Gn43Syk87KcVkS
p1qt95+Ap5lRVOCLbuwtzR6sn5QwtOes2eWE+/nZ6CAJmFjtoZdA/0m1Xf+45/1pWImo4IrdCFHe
TbXydpW8HkDRTAo65H1YU3Ksd1lwYcN5nej8GA+C4HH9PM5/haaL5Fy5dck3fYt1l0UnD9UqtXeL
1r6I8gkWEFqgOi7DRWX+k9jfPZVr2DhhX0c/vsHDvsv4QkiazGARxNI3sZgFOfO4brskCZUEpVsG
Lb+aECIZlwsbX1Tlx58e1Wtb2uOmQO0FysdWVlhUNexWcOIr0O6g8fa2Mr1tUS43lVqPSCCNu/1U
p8TENNfxymETwc5aXbM3gdXuqmb9Ib3Jjei9uPiq7O7LGmPjmeC386NGYzDD/QKegKKgR6G1u2Lg
LaESWMvXqLlTQgkSM23EOJjF0NfbEXKaExCLvAoKKFVw+PzlBfZC4HbtQLSAn4aVWN1oIKg63mVN
XyjWGjc7l9igjxpSjsqwZ9GHR5XzN8owyhbgdXVehsLtJYyAiwhq0zX37DC6QiVkJhVij0UCnkgE
emVAOOELQeqd8F7mjQPSc3gRFKa5AqxsaiNzAjpA6UCb1XrYOHqgF/09ZNaGyKbJ6u/Q8+vzrR0h
GAmx2e4lO7A130rpMzfTV6KluPR18ca4x4NHb5H3hHsV7Cki0SjLaI6ZfOeUvtcW1B+t/nIU7K6b
gvWctbZYp7XUAt/P01ol9w0GI2J/xbfD89G0bJOU/mlG8S1Tj0SL2NtBqVeDabxpYXC4iaJAnOxK
3KJ9S2pm/rsiqyZI96Fo/osVELzOPUvjpZM5ulfdIJLM2yaB/lMoRoKeoIkvxdF26QvAFR6fqPLW
LAkvKu+TyQU/H8mDaLstzvojqffmGEa3VHZZYrBUzkfCOTHm3V5hmEt0wKipDEMlSqtw4eepZhDt
YN/LsgOaDsEtmvBCjPQ7F75uiFvhu4pAI2miWxNMCoPqm6vFZ0J/j8qCtYykQvTCp2iKBLW+SifJ
g3O1Hhj0Sc8zEl/2/11p2E22MG8p0aldwR11vlDZiH7qG327DSEC1n+h4gSkf7ZR7H8xm/G15aZg
nQdn8J82ZlN/vEd+df/HIvAiFFS73P0vFVca9Xtz3dNbOlSUGz6EIIT9qSgzlSA3498CLTjClYKq
YywvvJPnhv6uy8JS5C/PJzvFu++UCGQN1dH0aqpLs5Z4gM130imSAbFAkkj7tQN+IlwX5c49DVcA
Y4b2dKHpDK9qQyydqxrHwzM82MhdN2lOAkV+6bYPSBz1lFOGdaeoCiZ/QdimfkjJ01VyrP0ASuGW
wwHji4PuAtGLl53FomsVSq3U3IeUtkBY9Bx+L9fCTNCjGlOliL7eg6m3xf8CN8010gukDtLlZN1a
fXuWvqp6AaaDp9sarZEVitV0e5y8dm27xeP1RmCJuha2vNZzevzS137vag3888JHYUbTDfYU4jBh
QR1tk6uV2kjkjBq5TI2CttygZHpGckRyfMKzWgoO4J0rn+6Bw7ggvrHRUtrOvWyIBM9JUodTJbNi
jAzqRK9526Lc6pRVWMbed0FrRNPcgESQeq64eOZWQox0ebAWPvGvTXFx5az2xBjmcMm3S94CVukc
ALbyI0FtuQDlWo83XGo/AvTcViYeG010z58huqhajhTNvOV++AeaJRDGV1NQGcDZjPPmzd5dwGXC
AUPauEikrBaS7boxm2SymTpcpOmkiCmftIxQnPJ4VLu2+yZbZr7u/JxMIYh+P642fZB3LJW0H1/F
7GSriGqOPktM5jMnxQmo3vJgzlsMeaVYWrjQkjE7dgo3ZHlNVofALJwSiqHH0kmrtopbWkzxxOSy
4WXF25nPcetlhWdsNEYEVH8ycs9//Vh9x5xLaBnCLuKSHiCVt3EAYZTOVKZ9jKmbB2qtfxOR5tab
rRGqEss33tnm23YcOV1ZZ1DCwqO9NxjsqwIC6MEm1wX8bVZANVTu44IAVTS3ssgl8dJmzyC8T6gq
uv1Si0HwzLAcHn0Ki5qX+dmc/j5wQy55nsisJRFNrTec8XhQsJCgbgzAzMIZU87YkDyPv4gfdZsw
KPq8G+jNuCsTSeHD2EBeU75Ste0DtzXACFnPgtQLaW0XBdWu+t1YMa/Fs9jX3g42BmgBpxNcNaeF
2/+p+hwH7RmkgrP5O7o3Wsyv0jY+KNnPHuuVx2FlDoKMBlsyp8rEyTm2HMMfhhStTdcbambV1VfY
5AN8SdzwuvAVHuM+AOmhzKzftlhW4HMO2CjU2GicclvktMX5nejebl9j0+s4LRmYCBuHloYhFVAX
3ZbwOb85zHS0iZsW+NEQe1v/RaSNech+RJ6R7z6LQeqX6tTPn61XT8hHJG9grbIiCXLfcdx9cVgy
PNlqz+LAjAzGxeVKIxu/hnrMsiSjLCKmISG85LsSFU2VpUrYtK0wOOjpP/63y7VPPO8fU3QHKuFZ
wZ0os3C9keMbkO220Z/gj9DXafWIB3D53yJgbIXTPzcJaR+tHJCWFy8GLqOtvp1owitKMH3WtoZi
FJS5k5D3JBrSeJWuyzj1kkXlmOHQTy7cDOzZpDtNq45MtecfSuO9QwBRWOcRtFw4V1a+dTiPPPUP
lyCusKEJi8q6pWReBMLAYVswioEd0E11sZdxmxP0WY5NiU1lIxNpV3AwPMimK3Zucrkkfrf/PSvA
ZYhEJWWiorcpcxcFsF3HrKQ5SNJWfEhsq/z2A+4g3kiI1BvRK+LR4DDRF9WxfQPfkwq8ouz3n5PH
R2DTS/K1VC7mvPdgf4B/RXdkI94gmpT9l2A7hOtd9dSdm9wjC37CyXK2zjCJ64Zd83SpXzKxO6dA
+MGWxTyve1zkyVPAeLnuHFFG9k0bg/YayxIandd9JlwBWC+4dUJ7VzsX2DqKP83XN8gqtQ1G7giy
M7m3lG8PuhRkTo0bS+Gg6K934KWZb5SLngVYeK01whV5S4SEPDM5D3saH+C2GhVdRxXNmrGHwnX/
Uio8SaxUyMVFNTnY8rl04Nc/PZ9MQGJNncR0N1HfsbzxJfBjGS5K7Xu11l/XpTbRg2DcPvqRFR1S
+Ad0wmb66mahYo0QZvp4rTIr79GpqJlh/WWSt0ClMdy5Y9xYR5MeK2zuf6PJFCFYVBRF7a/3oJNi
c1w5Au1KNOdTghDbS4nrLq7QQMoG6QyYYuUA9xJ8OcExOvvbu6xAhaCEo4jxuyYB8eTGtHnHSfVJ
hnrUme6o9Y1RERNhJD/WWZgeDgMmkImdeQbb1zgTbhyUXo1RqZ+mD3IXnwG7mc4hzOZ5Ey3zH+fr
advsOgSDDqHRu4jNvQ6WG7vW0NnETSGKVm+66DYun8YXBFRZfBy9bSeX154QeHomjiPQDFW/khNm
zTyvX6l8mEodwkVNp1exJ9v28ZJ/wv9gnuxOGSIB/szm3BLEm9MdiR2zxbANYI6UMGmVuCGyCNiu
syPBit/KfNfPQK2iXySmSqvrNZ4a79kqnhVnUIppA/Bu84xVuJUjbyVLZkJEmJDBcWQNn1knI/23
274w8Tu7DD3IB9pmG/OOrH8Hv54IxyBmFuGlKE3u5tQX0ANDGvaLr7EqrHxArmsGE5+kFt+8VylJ
IhqOWIUaUzeDohIDx15nZ7i7Gq7aF03KpyoGLT76GZpL/WyxW8WOdes+QfoRN37q32VrCkpfU5tL
E/Q7Tu2888GiXnWHcKdCZ53/+vWAi4LUMes6f2FirjkjPVSkxw3M1LE+asRtWsBOLGQPrwDUacG/
YLs8IkBXtu9fy1/eGrilr+v5+/Y+DLmcfvNPmU3IqXZ8o8ZmTbFRUn3zIPTGfRRy2+/aKIqoR/dm
CRRv1yYJFhnXbQVMG4eGBAGmjIsyaCePdJkRlZtRKFyemjp5V/BGni5cGYLQPcQGYcmpi2OZ+P5x
potE2E8XPT/K0BwHGjVVJu2hUaH4I/dWPTzXtl+TX1DM/R4shA44aM7PhGUYQum6/0mh1wbIuTwC
9QUasbzhrqJGVTeqY6x6CsCBfUG8oLPjDhOBrQL/M3p0XgFekeTlJrtD8uR8qWs1n3YQOaHTA+kE
BihBqdMYMZjXK+4aEIy93W+qREok0j65oQE4DqSmBEfwP5CDx7EHl3xjaTWJtpxmWTcmN0UulVN5
cblrc0Cis8WuNCecManbiouXpQMboXc2b0BjxvSS4TPr/m4xCKZQO0ABVJ1OAiO4gtUKWpARYwws
fa/fEZqZg48JHEO0VlTU5dXKFXsxkEDHYtvkzBGg1DxZCd8ahw+VW6NhYjwbm72dm7LouQge5cQS
tJ6yARPnqyjeQ/9en+w9sFu6YffKifYCml6jVmMb2Hm1BBl/IFOL+9RUYR7hMSwzwGfbnYwgTuQ8
8LQmzvDhTT8HDZRQ7eUcyaBKC/7eYoXU2eCC7Zn2kICKl/aTP+jpGyWeMZkBctN/8MmMIhOVyVCT
o9Dn2c0Nx1/j/hJRzBDaWmXMs0n/byXJqklDM8nn7LNPas7gg5HYZlDQvyNg5VdIEaPhWA6WRSi0
d0MXW7bgCcXz1nVESwJxWPMhzTNqEGNF3bABn0YUeopeW7VFKEVZt5HDTwNLA7DI5GFDKkGdHWHO
vyAQfOaZHqoaeMXKisq2yThceVg6+uKxteiRZJ6f67s6uB18dHz9fDuPxlNxHokWcXB+s6jpJFT9
tokrmbWBWpgSG8wXo9g08QWQ3vNOfmVNN5m3GW6iraFo8XQThY0j6dA31nyFQ1NytPWmJNqdXH4c
FVyO6apZlDr7nAZemgWGe6uHA3iy1udsg8zI2HgTb+QOyBkwIINXA5PX4FiDSyyZwGcQkU5iJ3QO
W6VVMJWg9nski0XrRCNabliRDwhz3DT61dyuXDnpE/KB+mv7JF6NDnAQjeF8G57UgWfthnAMMrnW
RGdIbKVtQrsgSRtf8gXWVIFyJk70NinTNcMmvBmM6OQKZKf6GBZ8JgDxiyeRsKLILGGdGxhkqJSv
ffBXkVkMHZmQkPtZTkkp6td8IcVmM/pvV3kZoPuDy832gkYwkQ6xqkZSKsFc2TrJC4YPhSAJ4+0n
8pHNZJ06oiu7YC6MnNca3GILrJISPxnXYMgDR1lt+6bngSTv3NabuI49ILoaWlOYHWer5BD5Snzl
0sdvtwZPU72FjqH3D04ChOhsTvw5hrT8+ATYdksTzBkAl7TxVxNLTM8FgAn5dzdL4vwZUJ+FYzVP
aKc60TBOvR7dFr4jS/MiY7dX/Iidw2BYHl+YMIKAiSmGumXLEcD8KziPkiY4vbjtk2g6Fq9BZZ+K
hKU3hsaK1GmquPj9beRtoBRqttIaUsVRYLTnZ2ntD87x7TE66x3rjGHphg2VjAUI1or026SSyzzP
8JBeFrcPpZVeuZac+xZlMnYO0uLOsCh36bYwDKMjIkjG4h3rL4N4gYFUcbNyq6oYFzCisPpNE6wd
uJRdUj2GZYm85bOKzBjd+Nwqhma1ZxpkvQKhHnKa9ggVILIL9tlOXk5CqrvgM4mtlyqn5aZzNMhX
X2wx8ERzEgUn2yBR49kIh9YGx2jX/8Oi/8nAanMXRez5SEArtFrg3TB9c2dbMbfhQnLOiSs+zfix
ieyDdSPf9SjS4q6oegvVyftuXhsgCKcClzYDbaZ9PAVSIPGJ+e4t+Ce42peN43wsExJRaZ0e49+Y
mP5A1rU8QUbEqWYpeOM/07Wgkd7TgUZXRDVjuLKljIGBVlcjbM7mBclpww6GnxRTCF8NBAcXyWM4
+R1zMRRH3bWBHOA5/tGVUz04lzzU7CyM4Aod4bUyp8cXZYkev5cv9hJp4xzNnMVZ7EAnlKjl1aX7
FloKWSoBNcCi+y1CByAFmXTOrfwaQbaKYnO1G26RwD1POk+BdJA+JxNR4E7QsKDM9nAUcNib5P49
DXBlJ+sO4c/uT1SER+B2pFA3FGFq+eyLdzOOqgOaqtAzibvrJKnf5gvc28ZcfDAEA0SAYAlAf3GM
U3UZfTv7aY9f/uxvDWuyPTVPH6enyU+er4qeExQQqUacdp2g8xFtnsi7fkX3bDNQthxILfXNl67M
rFjNQmKdg32QpjLfQaWM38EueX2vogEy7LfA3AiolNKlLNB7lkf9Q6tYB3cTqVGjHMqzH2JqeUfP
JFQxh7oAnzwXhKR0Ipwq+0Wztjo0zEXQ7+nQ+8rdvQLnwSwib/1UhX+sLdHBXk+M2xh3R/e0XSWJ
DF4pLwJ2m5ADpic+ch6ZEDS0q+fUhsYchzADCm+/t0KS+UG07sA4UOYq8O8dFREzfcDBGZqOCiC6
qWXs2sZ43vDG3a/M44RjfXQEJjy3Ou6+0/8VvOzKyDiupER4KSpaqlzaL3Hw27/sjm1vXsE1OXYu
MbzsFNS9vbkxbzos5ZYiKU9LupFCdepOJZtRF27gIU9HSCiDAe1cmq2zkhVminPhe+0Vey42SPza
6z8KabYz/ImI8wactJm9GwIYe5T9qrE6iuT5NTDaBaEo6A6yac3Z8hEyffRAtudw4IHR4iVfXfKu
doTRyKpSH0q8SxWuYovilDxI07Ij/HYZVk17xGHrtD9XiacxiSFowMa+EAzDKHE9kPFmYQtVuBrE
EfjnFxtzIlQO5KsOvhFkrZRqPrRTHTys1l9ktvPUQal6TllIMS6GQIRs8C1xaAIpRfJtMNjUjO+6
HHB6jhQkAHB015TB4IfZuwGinuHsqVTBGQI6JC3/Kvr5bNTr2QGktnE596dqfPJBpA5GhEhgXgjG
x56tdZFrNiBNMHOhiX1PwLGA19MbhnGWmiZHWRfacrTK0m9QoEKAooQOi4W/WjHvNszDO4Ng8Y0Z
3zVxHpAYMsLOP7SbC+r43fiY8NTBkDwE0RDyCi9XnX3iFQCztXSWOEyrLn/wIBbnzKOdaoKO01Pv
ULXUGowAYASRLsft8YxA0tS+73ApyCnzTWFAfvO6GLI5kPRxZdLlpa/a2ta0k5jUD7dwIJpvShwd
0yzt8M4Am+p1iVpqrLzAMEdOrGNJiIIpvG7Byi6K/LKfVkfjsfotXk3LV0iVNUeRqJHESaoBJBJU
2NmQ0qT91EOXEo0fOzvqtFXVsoI6EXNYS+3BuomYMtXEQ67Brw6PSqy+h9hzYZY4npzhATfMQqyR
o2lXXWIHugVF/kwz2wuAvDl/gVS+t/4BgK+sJt5qekfLcimDpleoCSOSIfPUERTDAxN+zRMSUil2
DaX8CIU6IDR885W1q4uTT74qIAWUo3czfJ/ku/1RExk/MFxJxu5mEnXmEDJS9X6n9XymtCsTpw3D
80VFtkbm8RPbblhQ9MKl1V69hCTwWKFiba7C0kgYw9tndIN89OBi3BnXCVqxUrb6pnn59YQi61yd
a8VqVGuxHZd8x2++701f7BBQ3Tc6h7RhbpS1qHoF+cz+xztGI1X6inerJuIvL4tAgZ9dWiJwnoyN
hOThm/he1Q+l3FWtV2QqIeiOtAfR7xsZrgrnpvQE7rGxypqBw6YSigy1BeaRir3LejGr+4/SX6eO
YcKQbuHTsw1JTYQ7BbXIBNDHE/2ksTd88K8Fh1RPyy/huP/ewFsNk4SLJwMmpha67HEICwuypVGK
RdjmDWf98z2ZFWXszYZ/moenvk9MBSsJHFDMxc5aTrnFAo2ooVor7GoXFeY8omTC48KzHusKdtkm
JgbhfrTVvxyeipPslKwVd+B3buPwwMFwHrqJcRI+e1WqbnJHC+MnNc/KV22Pr+cmTpORSU4sfdW9
R1RtaGUKAizNkrz5EbIHBiocNjzWuzX8sxayn6lrLdLbdVYJ5CZ+6pbZtK2KfQm+vo6i4prCC/DG
Kg/tZNdRguzoXYzYzL+im493W8pbF1sKXlS1Y0xcKvLMgEw36IYw2xtNuGRawI9sufi5UF3MjYPp
7BxozS8CQmEKuVTWgBVxfVowiWw6jnXe/VAWgJ0M5BRI7QUT7baphxVfXCMQSKdUOKAvt+SkiOFk
QRvN0k5ACajLnh+mdcoVVEsjWS1R2msLCdnzjUO6y1Mx0GkDCgTxZq/p47KkbWk4nHC+XqEsnVl3
u/7pBmnoDkz4DCAhEpl+6AsX4t2Agyox/rQeTt/au5ahUA2j/GYW76CGJW1fhtHzSxDLB/KmvNvc
hghO65fZwq/yxsQf/RGcU3ePnYzx4UyhqqmgzwFRvHNVFZ5ECEfyT8vV+PpJHmfC84N8OZKfyvDb
+GQ/sd+lWIFSXa8TktAeOPUZCJFr5x2VJtmdx3HaNcioPNC4ukecr+2HpMW8c3402FyU6D75N6pV
LeXznEedygsig38oy+s93tR6iNTtnWhLnjkSPmEiSu0/LsbepM9rxA/204im5cy9p0/AspExxt+K
RFCerCXRNzTAkTHyQpboQCtzdWRNkL0a8xoWJncCf3LgEWnNiXcYm0xRE2rV7fKPoYjIBKQ5/VuQ
zmn2ARcibmihsx+67+n6mP3gupaSNYnvnu5fxiU5Jv+58J4KCthtl0scd4SVb6r7uEvi3/BV6nmz
IMNN3HRfAwp1sKgTL9xfPAsDSf87DavVXz6qTl9F2aaMA0wk7ov55uWkYfK+rzlUI79uuGeUNz4a
3LHD7rWePR9Chc1duS4QWG13xzvnC12wfman50qovX7wheG2W9HEnZYm9tCbFARnJ7bp21i+rogW
QoTZVMImf0dFZJu6yCptrZFP4iccqEshLzoNdEQozIA+8qQ1QF284EIkNMaxD53QAFaGypZ+5+mE
NVFKjFG8aXvNsw5cTaeYZcEg0u4+R06FVQd5PXx+9xS4ozSh+bSGE9AmUrguE0k7wR0ZqlRTFzti
lpcyYxZcfHXNPqucKTCBvDyhr8UpaAzf5OGp5Gq+CvEs5v6m8rvuPvspxz1hhINAaXvOcQ34SzMr
cpArVHJ/+/IQG2rz90BHXFPtXob8AUiNrbIOj4yW7FUGSP17E4YixJoZl3OoFK+i8sRu0dM7ZITo
1KSTLpW5FwLu95xNp4hZjPmsEPIqsHbJEsGqAcu8aUamzgHsHKBleCGeD/MbhlceazJV8lIprGNS
wG6AcjNQvhyDlXMhhr5oBg/JW2rt5lKju+rRfwzcsnMCRr2pPA2HLj1rA4JFPNxk53/Nsn/nOUE7
OIRupL8GX+ZZdoa6yl0hY5JNJb7Qf55bGbT2Fd75y08EvlwkvGbxGuuEIFkCdgGDqpmEMVjwVmM2
dqckN9EvYO9DW+oLfLhXl4jNqhKD0tu535gRoZ2SOjnyMEzmPlt8wg+hGh0qdNb+vY3lbnlcMP4G
9l/1FVu94JQ4uNb48323Fa/cXv7iW7nqz8OeI0sOLqGzNqKsWPV31mRf5Vm9bv+lelKBychYcbjT
JJIxE77QQ0Kz5bO3ZCIPbhi4n0G+MkLrghlUN1pZdEfqOVhP41jFlNpH7mxxVVaxk/dF3hChQSnG
b5pkM60uCAmv29ts5HHBSCUdDuWY7JKIB60G1OtyNe6UOx170mYSfQy26TwZOOYZpqLAk4gj83VV
JxNJjLmNrXvvoDJjJwJzmm+du9eaN0tRN91l/ClXgGdYufG2gwi1YMlKBQHLESBkYShVVF+jURXQ
Rd0YNFpQB6bDfBMIaPlvVPCiXk1+MitoAAZTWvlxYlK2YfYRBa3NNbPcSoz8D14kOi044zWzm4Ki
dUXFunUnO7U4ax2SZYv/Dci640i6M890s+YgnDsL7a51iCPcWcGsXZpK6knxOUE6RJ0xC6X29v8M
GU1L9rUT7jITnKG+bRglKJfACDjPCFoCKVKlKV8/BEs+uzeSFY3u7PXI/YBJ9KyCdkvdqZ6ZAC2Y
ztFPEHWKlvFk/Jq/5CZiht0qCBZ0OkLuHwprZRVBw6GHsJQkKg69lQdETgsT5tv/3oFgEg26s8N8
7AUGa4skaJfGLDQRygGAxJmfb0hDPphEOWHdKWgEdKvWrE9k5k1Ab7QyrMQx6PK9DZ8ayYTV24vD
CDsRdm2lkFVlQOeypQW2O2FN/beQF8gb8CwRoCCSQe1H78yEJYmzJvEKbLtkeZpYrkwgEBDAPInV
WcbDlzRK4D48GO3sa2NYPZ3IaOsmCwuYi83lWBZ87ZLSNayko93YMtBcKd5vED0VHoSz44goSpWv
sBcitQDUMvYYYF8FmC9HrrBicM/Jz6npNEr09D2ZN+eNmRqylqtl2SYplmgL3CkHdzZOL/nKgNVJ
nYC0gVFzSag8Wqk2TLEjr1FfzuY0HkIhlZKXs0mnYSo0BC3JFGrp+ckBMobWf3WdVxQLvaUIlspD
gPSokRLwQjXmqr4TxF5T70wmBgni+k54a9z/A5xx4oazepDiKXFHsGM2Vq3s3jBeq4fBlzrJOTtd
TmyOxjLq+vnZWOUe0KcgI9aUagJvF94AcCKGbAd/ocnIeyFfGYULfo6MsYib5zdG9SGGIZD6yIWp
d+a1WkIdEigFrpBFdOen2r6EP1u2FWjawk69oKks15Wqpo3Mc/KEiDlCgp2Y76DuRIxkMMkKgEEw
OW91dv/WY0yO18hKOFnZbZnijG1n8OkqPm2GZTo2U2pDtITCy5RzmOqRnQmMPllW2Qaks4bTl7Ss
QUMnJU6GLkTj5Di5IIOJPm1iEM60v4dCB5s6K/qCfP8I5Yc2nC/alU72j3OlmaCg+Ds8xXJjX8Mf
SIGJQ7ZyVTiBNgTuxbHlCR0o376W7s7/THknZA0zIbdCq/nSsqzNtu8uoHcCeZbRiv6tjxDHkIN2
sxadaMTFY1wdHsBRran8vJb9mGn4tL+hzAvQ0dELifxT/enWk55/g0EXy+yA6J2RAkxJO8r2ab0w
/fe4edq7V0WryNSdyWx7y4JP94FCVrFf4eaUeuNTj8i1uTfvBdA3e/OmGhlhXFH14go7ocEvo4hm
Cl4kGY5XsxvEUn+ubwpHPITtS23+9bbUBntI/fGG0t19g5tT5Am/tZfgomJwdGb42LkfVVK2Ztmn
Ty51TZ1gOM+23QTLm3EPS97zwl/5n+gfUMCCcP/Au1NLPPbz7tQE7y8qL9fuBQxKehJyN5tcHkdb
TEWQP3b4qWyHKL6B2TL2lzR3+HKd/E7Gh547kZvxtC+MjSjvSnQ9oqdTa/iWyR3xqlOds/Ldi0Ex
5C7ZQxIYNIJ9HYBcNohSelFoWzlJq+d5sP7m0XX9U3HRMyNmhwP/MWlmf8w3R5rD5U64J3bjFOJp
5pqL6ZlI7MLbvgxU9E9BbPNTs3oKzk7yIuVXXP25NfvYiWk9LNL1NikO2x6opC+lRMza7C9AIDtm
KTby4jcNPy/TvBqZW8JbHY+tYX8GnxzvKb54jrg2Dm7nScTtO0HkesNvavpOMYVf/Wkt1JR0vs49
VOxrTKlieFbUET4zyTZYyE/rQ/O8RV024YjswkzVlIrm0z5Jo1Y2aanLwTx5593wyRa/U5PkKdOm
nDoqL6xPpr7/1lnoUJ8bMJQNMIh6wpjACA87pA1K65v4uDkmDQxK1WISmsltKnFXZaQo8JxX03YY
VsSG+Twp3rCJyipA5ImFEa2F+xy6o7pjBmV8YuKOPkZBwCJ9iDOIrF8B+pLORe0Htcu/0UVxX7CG
ryAyptcMTIqA2mg8/LYrW39GPlYl+ixh98TAsYk/qg9UgqsFn6kPUSP5yezvDcFYencPK5gahQuQ
OGcyt2IvNZ4JUtU5bCKU/GM833+ciqO6M+5F38m9nDpQqWEvEq3ZigTXIsh7xS8v/Ck8/5rg4b6I
P6ZH3vYtdel4SrfeAe6S4Wvyyho8/tcbFVHkJHdQ6eVAdFTRv6QmA9cF3C9Gt2F75tgphoRF8Oq2
HKa1mZqo5f1HIwTDKqA41TbFQMgpqb0zSI4nbG1VGLWWSzqvykNv0+bPdLgNv6S4sk8mn6gtcoHi
7fdqbd4NGj5yI2snCUVAuXnk1QiYJpQ92189Aws5TitaL/wZ/vNdO4duNiBN9p/Y1NclEVGN+O7u
mul0VR0/53E4/pva2ryQ7aVhZGA4vsc/gj788hQU3dTTdjBXTEzs21CsaSfmVnoI+dX/m5nXLDut
lne/nKxNWQTfJxc3Xa2eR9CKgp8Maucv3MgWDEANzVJ9rSy5B6aZf3qy16Qy+2DMbDTN9/qYzl4V
dw7dVpqGgHuUvBiVQfmL+/IbLTBVQTE1RZ5B/PCk1IBFZumI8RTcbJ9fl6ccd73RVsMUPkUqcxFS
eRTqZnQm6ZJ+C+mJba2oaruEFymg26Y4Zag1nVcZlqs5sWts+iRVd9cb5WX37BNGZaOdDe/30eHv
Rpe404uFkyi+thpeqRTdKT1CndH6AXrrUCxAaCI17y0PcoS/NUcYLGwsAg7pcQ2QF7jTa1C1zo8c
3hXRFQotvrim9pmTXn1vgOgh2RRQX470bOaHR7xL7Bgl3fAOPd4twwqje1nOKwtxA8i/V7H/RpJA
vi5jLsDFWsYHDN2KqXcMMg12CDyxcNrh8HRGv6KPJ9IFUdgi/DyCNY62O7nfe1k7fySccS7yDrfk
gDM7pvDkJ14WCouIFknxW4d+kNG6ZPIx+8fuZj10nAWU0d6HbnTWMX69sifwncsAlYBrCWAAUB+e
/0MpS1b9KOTQ73Ba16gqXLOAJN1bX0v62OYJpImSULkFAbEDWGeljh0IcnUVC78PgI5cBop3ZwN5
Lv5bTFygL5Y5pLkpR3LqU6MjLCnlzgPGqHVgjAfHDuHVyPhJKXldhaUouLJwaXPdVRv02/hU6JHF
1zHBMD7r7deKmeVmUFMpmTLWDnhrOCH6KEsgsx09i/FbwBDId76niTwRboKZo+X/Mk3RA/hs43a4
VyC8hDVdh2R3VaAchJiw6nsFgZleOzKXhqsv5hSOumDmJsh6cbCSJC7GOGfYUIuCx+TfOH9ITOOr
2ry7gYsSHEaH8pn5qWLn8Kolkhb6Ph02ZGB1HHoALbQwJb3Cs7tbTwHWceTqlr4/jcerUUqi+I91
/hqdT8CRFP2IJgwKQp76e9dTviz4KVoqhjbwp5J8raXweW2ngXh9Twl66leBE/NROozjeefu7qBv
crJnQlVO6/vrw3Z6KqRyDAbP0iDl1hx+AFsQxAlGwsSg1BunpFWMF3S6xeL9NGfHRfumiYstAjHn
nk3JsMhCns2jVMekGYeEU9SYUrcq7inryp3JZInApP7keTecA8NmKdTUpJVupnZLm+uSZPiC+cdM
/08CJ+DK8tWBKOTZIQAfM8eQKPkPLVL9wG9KutRV1gzNBUIp64o5TfF+pPwwPeo327QXewO4JAUE
51wXGfclY/hrsxsze2PtRIpm/91qFoCtZYV2YQWPXY5kRCOSL1QDLmKcWnRh/p0BVwdQq7aK/V2J
R1Mblxrs79PVFSYYdhnXqRCQT8G37LPGBr+icdiGx6oEiZnUWJGG3OKNEUga+p4j4WPbWm2SJl1L
UVllhCSiRg+s5nziFpHxqdfPirHYU2DtZLSfxMdfM6RJ6oxAz3n54Ibi3rfi8MLXL8pnMwXwt2+V
6I4uYSSqsqSZKZ/Y82Us90JoFxAUuF6WI+z9MKBj6njx4qyCCfae69KAkbJSPEjDcHvru7scddRq
Az0zURdLBaPcqipgec2Oe1ahp3jfcBdmM4TciW/C/O9Tf3XciGpSb9mb6NlCWcL4nNXIG18G3DS0
5mYczlC7U9n/SZYfWaZNlk/g1FJZxT8fWJQ1I8LT5rU1lVq1YJr9j+BLSRTNqcr52Z4PRtUsh2rI
uBQe9YTdVbcbuLn/1J3qGAUGlSb4nPTxpZBpn+AdIR0OZi9cWhBuNguYOIIfcjCtr9r+6lQVIkR+
1WWwagBmGm0AuKivzoMZdThJMhUZ0BLmUgGrIMfBD/etlasxmXIxsChF0YFe72L0GRa2e3hdDAYP
5iJZBp8R7dWL0dDED0CaJmn17M8m/ZIM3aoerewEoydxmgXsnZvmCAAdndoV3eBwJfP8ke7QjHGR
4/WeMcsnqUHS3TbyCur2Z3f+zm4lnP/Mz5pmJ1zagymGWghG4HkSHCtB+AaG/Xt25QQVzbRp7phJ
MmJa/Bt5akJzAgm7P82mzKU12D7V3SpBPTp1VFF6rOHw89s0bQgrTTrTnIwP4xgDTUYrUvEPL2OZ
U/pVS6t/2hg2A0RO1UBwaNjpilBgocY9JDNaJqiDBkAdipBZKpO+2mhLjobdJ/hLUalHu+lgbY28
ZAR3IDnfyL97blfpKHCKFZHh95OAXP74TYHimpr3wUxTPmG4JdhDvx4JfxD1dC4R9dgDJZdT4Yap
mNcgzoJQ5O0NeTxJE3npMGdDqR/R0XVJ9x9kvX/tj9anqQVFCtuwH79CMKg7VY/KbXLSpsQictgG
moSg1y0fzI9YUo3sXrWdDIxpJItGF+/3xylL7oj10IQg2BvD1Z6R3k3T5e8TYvwcx+4jG0HGcLTZ
4JhRvod1yvvvI1R1rJdNlQLnB99Ho9lJ9QSXQN7ALtnYI+pSCEemNWgHi7tK3Ms3amvuB21QR1R5
aWSb+6n0NQcBWuwNAm/QSeuQfn3Mjer4Zi/o00h35IYrgUf8gfEctIc6APsP69uBoSmLyAhLwCyp
ADHBgFQvVRjQEd+PLsIfAc4bc/HfUXYX3hLLcogUkl4s5vEVzVmKAzeSBEXyE9xxgMc8JgPbVcqw
BR9No5pcUO7b6DBwJEspCYJwMT8QVUYtyEZpsi3currno3KB/4zRPSMR1xSrS/BKGgwyQr3TliB8
R6KNGy6U48gLaELFc31DONou663TH3GCdNLZQtJRXlkHquIeGsA/noxwMAX45wpAG1JzxEJnDaE8
BvkwuAJdkbYg98LsglnB8NaLnDuUy2t5YyMTt2La2opVmAEBxhwXRsvASMF9jTin9qbNBUjx9j9o
Tz872ES1ZUnGf7zjMQnvbfk12GW/eh8b7P3jK1/IC8Bq6XQkURYI2NyH3UxBsRt+bMDJ2X37l2T3
WDOfCH8HrLqJXPFahLv2PtMPYLfNb2zyZ+3QsgO2il5dDydNXYELUXgmUv3B2i3/NS7onY4mpKcZ
wDPj6MVW00LtDCzBLzcGWWFfgznlxC1FR8+ubessn5gf8RJx9JLd0lyZ9bst4qDGGKE74k/GkV/+
avr+sdyQnx0TgKNzJ//8h2fxgrLOUirNjuAxyo6E0lorid/CpN56/Xu+roGjfrvzn0Zbk+jn7dUv
rmGSa1cd3jdG1yCpVKUI2UE1yHwtT5Ge2lXweOmB/fsmociNbobawzTYvMTUQA6pKiFtv8U7oiCF
56yg+tAtK3h3IsWbCrJou/6+5sD6PiTQbU3STbenT92LEP0yJe43Tqf6mKx2se4+A9oBMs6xTZIU
4lebrF+bWv5e+vgOkwv5AVLsUxjLua9mhbkDz+7cKA7H6POWlpDmHcH94aIOVQUOimwKi//mal/U
ds3xXjC3urSxG1paLEBXhDhna0FR/s3I7k6tgVfhNnp+Wx1yVzqzAnwgyjEJqYG9UOVLrZkRj1LP
R9SAeT0652sfBxY6MqUkON/QmZ112mDEc/9VRnMzDyj3AoeSIYz/WMTSmtk0VI4Jkpk2Wgp4xqCB
AK6hnfdk+0KoR6/AM8nUc/z7/R/SqSqvPRcS0HbQTkOIyZIkcAkXgtz+qi+XNcu8c8m4Y/exflms
aLZqoqLIEDBnUAIvmWSN1jaCbVCkvLDMkLAUpR7RZoABP6plidrRONeM+u+afKf0KsU34ogHcB1Q
ePQ3GTmUZmMLtXRxi2OWRWFVQrwLvJ/x3MPwY0rb+yNWC653GE2qd1/plUvWNDTWzGVBUqf6d0zA
4n8E8phtLkUyhxa0l2e9NRmtgbt8A6bRAmROZ3jOCvxB6hUY3CYrfGK8s6O5gACiH6sXtzOl2u7o
+TmYzRiRUHAWcfScdjZcgPLr7au8hIkCdwDW5nbdwlXA/ipyr5Bxutu7h2w7ZcQ26SHuel02oFn8
T8RCjZxFgjRYCHXTnSW9rbtgS1M3FEUmFe34Fu2+BfEbE7wl1RWfmztbs+PH6G1+kF4I3nE6DAcH
dLWj+QnERcktZgAQjMx21Knbd77+XdvHS49uVU9I3QCro4f3Y8mx3kMjqVtcmR1OplSmDkn9Gx/y
s7JmvCJsM5zClNgwKeflfRj9ZfAVhyo7iVYsIIx7X+2Okufty46fnZQLshajMJBG72dGJYRBJpHb
N5wBxPb6PqkN1VdIGuk/4nfsh5nPB6h2xt7hht/XATA+uQYpbPk6FB+Nte3562iapT02+Cr+rT0m
4QnzZw6pLw2MuYZvyaekJrtLlvNJ6DqNZROVFI4OPsAfEQKFeaJh29FNThJZSZm1zpfdhlrAjWXD
Wx2aIGwF80xnW47AeG5RRPqEx6bDYj0fON1uXLiuOUkyfd27K63m00LRm5Zc9wMODlmLgBCsrrz6
0/fc3B2dMVLDsyBEn0+f4ZdKfvaB6DOLFgYHcXXUodVninR7/KUH0O8Nw4coA3lA5KqdGljIeVt6
1HCogfKi1G+eeVn7QRzFE9OIcbgshAdh7B0c4VXMqIHkCP9L2+TW30IkmkLYYGEmBatYNWlW/JmA
aefII/JFFUo8lLvsSCyi3461W6RL59f16mZnT2OTKlHH6nz5MNy5tvAN+VGTAkqXHQMcIsnKNrxl
CxuFVTiKrQfQ9jwrVZZQv9mmC+cRiUp6ZkEHR3lfqK9Qx0xtM8XED8srlUjU8jISoEkqTyP57F0F
zxfE/DCwbJ5pQlbG6giDHyptHHu7BWtZm7Dkfb+aATrKz7IYljHrwRwsvlro3d37Ex9bDPtrbIsh
B+hHN58xkcqg7Tlpk0lQurCDEYyoClFUm0EVfTOs/+w02utVQKc58T8ANkdfzv52ywgTLNtN01Fe
SXRyDeISZu9c0t98Q/PTSBB+vcHE2iG8h+UaH6hs+6icSXZtV5J2ZXsEc9t2Swup+Ehn/fmJPbn0
cwV0ucKGOB1dl/i8eIb102F1n9jKhkyv1bDkSIH449IjrLihbkK+TZHlRoKLNllWY8dZkY2P9gCV
3Wj99DLngjYjHqDxHhjLRr6cnWCp+HSwNKASyJ4gYORoaqd4JgcMDXYqh4Ac/Bm2FCqQmQEg/cww
j7lkO/YaS1sB6KVf3mWbOM3GE1mqiD8QKKyj4O7jZtnLnCo45Qf+cjtSfhbtIAYKWI7Mt6Jyp1hc
1KzhrZMXDRAl5E1dza0FOZhRxcvCU3THnWfqbApm+4ymGAxEKDvbiPSNUKiwFOgOf4trlZP4Kfh4
k6PGx3h8FrIeKmGSaEzk5ojpnqCIYmD2eHs2gNJkcKSdr39poTcWUFUSwtWqBnhMqNLmdX0GMztq
5Ebqj6Re6uL33haibah8l0qsFssRwmgi9hBLwUy+IjhydEcy3NhoQ/3kivsNncx3SPbb2IjAbwqs
8rEnQqfTP/Vw3OstxKpIUsUKolM4G/FBwi+oH1ObjWKoMuT/yDP2Uz2ZBcwDywgSBDyxL6QZO0z7
O8f1z6fhmqExKpaIHSTV2JoW/MNXXLzX9H99rMx6jsLLABMhVTupzRnLGYTYYckDAkob6oFjKP0B
T25doo6rC3AEs/WA9SDembkHPC2XNslYKh0shPybpwjsL40IKbMCFbXSp/6HRw/Uyj527UhmTwfA
F1FJ/sYcH77+PUz+uKQUaTwfr+/K232xCUJ5pMyEL1T+F5fLJXN+CZTIXKG3Z5XJDzaOrGsRUtyX
quXxa190Cwlso1tXriGa3hNQ26Dz0ScMfJdKpve+Ihw/rvS0tUPZ6UtGChbiNvq01lmD1QDuBQI0
7vlFNswB0NsPICLUo559DOBJ21zWoJAfBOPSUfWTLosKZ+3ZgdqASRMnFyzx54qIoMRT5DQt9/UR
G6LmiqPTqi9rkQXJQBK/W8JaNuew3FiMFTp1kZHy3UBQ7h7mPzbT/DzEkfBcw1Lo+nZ93vSd4KRd
mNtNqKF90xmGVOpTdn5JdkwRF7UXvQFRuul3kOnIcVNyz3jjSAH6kvhr74RmoQ9069QSyRE1PRor
4HWF24sSR9RBczy5qpsJ8s0aikhXE0ZqVkVsQsD9UO9SszUK4bxouXWISfF6T6T3MUmnGBf94ExD
MwBAR9ldMEJizjkRrx7mMb9cQmfYijsw+eUuEDpKXiX4iezUkYBR62mVfmwK3SP0uiiP6q974GdU
6C5y8UuTz9X93Kp2q1KBCxLZcut0GWKF8QoqonsKpFQ31VBqj6Jc+2rx5frwg/qa0mwvE2DYamD/
rlnB0cjQQAzkOi/fBAmBEzwXoqFHAR5yCtIj9d/bv/gRgknqLYndJCfHWG1nyjpzrK4GJIXtxzwV
dhsE9ZxQ4l9hmnXFzfGXKVjB9SXMKUawuibDaEQzvkmONkXRAWOvI2FPhH/HqQlaMkgB/Miyp6h8
fjeP4nhHzrJt/S+8TSLw0fCp2kPkKVEHh5nwDvK3qtJSAUYFjlvavdbAnG+CSF1LFUgeKd7EZhB9
Gera5Lfe0FhEyjkiQqX1Do2urVTxOyh+s3NBMFtZiTMOO24uggBJIJNz9ewM0Bn1+ijk0hZGwVGL
g00fN7PG0OSfvlsf+iQZc0QJdFK35kkUlH5+l5EmifGpPXvahSctY5acvU4Of3Jp53aNu9/cbjM7
xjp2Z1BujnvO4Xp+/rL/Vm+8mJKUMm5ylTS4dNt+7I1zxc8pvX04P7P4oYRnZKUM4vme+Q7FOofD
1jXy0/J8cYJZPp4/v5rCBF4xGEtWJKvTom6XhR7CiCpPPn0rzI4eY5EQrp2i4E2he49gFJ0INxKZ
m9D3i8WKkvuYMstBxyjzl0EZ/syWHGTOEb6zjU64zRC3jwrbLtSPVaEiIbE8By8ekWDpTvbXTuVq
EOrfmoQWMEYX2hWT/YZkFnVmDNrAFM+MYFcyxbE7frp6Rq4rDi4uyYBOMv0tm7wotkGzDdzr/ssg
i+iKhoqryEtyReaijuig5/jT0okuIW1pSUbWeFso04S1grI1igOYAc8L4b9dXJvF0fZCr6x4WAsa
nIc5rFWYo0Q3Evjri1xbOpr7lvuYaZaxqvUGPUY7tT90SzqjcWEjJoTS5Kd1Y+1ya1ome2Ef/b9V
hDDw6pl/Srbyp0oqhij0wCBs5435GZyO8RZmC/BCxvG9xf3Cneo8u9ygrRDl6Ty4RKNrBcNqWIqa
USG3Csbgtft2XSqAnWTCTT6MCV0bJVslLB31797qV7XwCQVFYULv/V2ayfTwojb7+FXiKCX2D7SY
HoDSc+NhveMRFvmxm6SuBZ3zIy1Ke8PeJvdYPype4IVf0mpQvb8ZU80n6P5Dlu5fiSSe4Mu/6VCJ
/XlHElqttU2tdegVm3BxFRKPsfgqzauItgevB/bvrVmFNCrtHcGxGGNy0N4hsi51izh980vRbE+3
5BNH16vAhaHOdL/xd2sih+yeFAFtpjiFH8ppxL7IWU0VvlSQVKa1bil6xEPNW4OkWaJBWELjxd/3
hahzQ0XC/ix9N2OqYZbU72zjz8oiQN/gjW8bAjuSwctKeCIGZy6JLRTP+WmuKzrwOgfc7BMcBer7
8MQl4LIs/BCDKq43YnvwlbQN9t9VyX/vst+yQGWed0SO/0kZWeRcglodd13hBPoQHI9ruu4rUvhl
wiSw+hAhb+2rzcKy4EwRTq7z4LqmRUPjFG2NHU+iUpgyF4uwp78AEwsDH6EJO3Ups+L5VW4O3bkF
JLVWsm5TxQZb/J/wrN8jZfvDvARnm04i3CAZN8v5KndvtYfZnOmL2QRQiBacze6t8iWFgNxb8UWw
w0b+yukMas6Wm1yd7VlWAixv6Bk1yITuQg3FjzW2PUb3lB1g743BG6/D4Od9dIqggkKuVuQFYysl
oEFxo/lqzKs23xhJqDF//C6v2KISlT3qNlteyVwSDBbtRZ3jxDHK8yr/lVjm9NObV31r9zM9pZLf
NnuwydwQ07f4wI9eDfWZLuoc6gIoiEx//uEHw1MCua7j38HNfXJEOMCqKTEHXIj4C65DKtbvysPQ
J/qXzToCcizb3G7RniNktRpn9S4KkZily3zUOiVh5+y8424jH7lzaKfhX0jL3kfHYmqJxIJL3edj
uAYO9QxYT1pdxpsEiQBLslxZK5/ZEfah5OWsoe4YeKly+wAdYz67H0WwbD/2Z7w5QvtloT63tN6i
AiWS8i3X8pQbwwy1Kwg6sFnKZIfKNJ5TG531gQCF2khw0wQ9/K+kwH3e4inMuu6mUx1LjI2Vu5RY
t4it7ByUYUcVCsmwAl/UyqYrPpVRWpGVie2P/dTp9q4XWlSVEbEXIEGQ5gk7mxER9jMV1wJs41mC
ys45bYPS18IyDqQf0o7bJfdLXqS5rbtjDM5vH2AcbUj50BRrjpqPCFWeSeTcTVbJbNTAluF3UkU4
OWgN2/ufo70+sjXWjMyfO1Q/1sHUn6JCRAYXutNAGxaLBIM+zwGJ0fXpfa0wEay5zPqJs0ojxCJt
dKWG1eqzHwOcOladB6PoAnDboWSJ9ArEMB1AqfKC7bf9ZeecHGPB4qvn264bQ9YtKxMDZ6UWPrSz
PTrR4puEEdutVwowvzYyo7tdtiu8mg46GAsTBRzv11/iF3mo54Qmznv2KIquZjMbe/wchfUqX+YU
yLtLCKnFIteyGh28DQzyccox2pwZIq5x5U+Bf404iZl8n8nBWf0+21d/7K9iamwA17pjg9N0yFXX
2gghf2FrRWA9xRGIMioYvmv/R1CnYhBh0WQCAD2skxb5ViJE7xMWIbZMU0ZawaHKQx5JeyRpXsKO
yfnE1o1gYtW0BHbZuLVq7wXvTUP2qBBJR8/BG/BolxM9BIu4nE2+udUEmg63ROD/JiaAZ4jqbEJe
kUWceDyxLwEGJg2zGpYBvnv/XFNtSAyWODuZt9BOEqPo89ceNNLLKqLpBKbv9N1FLsQMhe6dtxG8
N29XbnpPM8Y45+MQq0hogijnflNPMqw2fpEsUuQijfJanVi6hOof3R1oeJs47dMJqf31ZGkhQxjH
uQpHGKNmSqFP40MOMOJw0QMO2J1cPHmV1ND8Al5ObbGGaTvfDjlJaCM7Oz+1IMnWKhV6ZkWfObZk
N7iY7vTDXmtrPRe94cD1QuAfk84xHg5qllDfTWvZM5dMUiSRgJ2FyNMcsUXJG7gKS8Nh9j/lm86+
pELzLa5wAEq14fQrfgHDgwB/7yPtTOBQmjidL+K0pcWsTAFSJuUsbJO1mZEx8DcSmAWV30ul7jnS
dolqeGuneiFZNhyOYG88L94yosPOepBfQD1ZYwKY3mmn/SVczKBP6ft6TeCKOKVMF3U69SmfoPft
3+za3gzvgLj/W/U7OL+zzCE/yGLDLUfLGDZCdoF/2nCtZmw5IE6JmDUDIMrsNg/NxwxqSfkFpwGc
DaM1H1b0d3ZNull99RquFe2oALNinWjJkJbxkvaY7NFR/v9CQ/o1IdzpMOupo+PyHU3TVqFOogWr
jEtuAfseWlZ017TR5JlpIpfvNnJYQE6Pgc4vb8L5VTnJWcpJDi62Hc/3kExaWE7P+4Cgu3S1bJZi
sr80gecegZVAWWsa/JG+I/B5yl1x8Udoo7jL3u3dgrGIrHYMy1uW2YZ1xOD92iJ1+VT8UnK6VXCG
SXTWN5diSYZvhNdqnSl8N5QVQdYDCagX8zEe70KMP5nTcJgZDM+8lQM5J2i6tFWyoFB9PNywMQab
GdR0MfxUFAiT3uKvgnK/8ASsDxcl+LdjI2bj1u8AO1CFf8KjmvxRHACmenNDngaY7t2AafOAOYNG
GqmZlWLDpDPgYtfvrw6gdN7cgaUqQOl5wMkhJyuRUVAQMG9JzTb23EoQHzANourqwghsseQ4t2zJ
CI66QHgWnpgjVmaiiX6fcM3/wByQwulbjvcQ072/1PIyWFqhoXmX9pKD4n9rjuS818nzTiygzATT
13rw0M++NNHVMLte2ufyB2e9W6uqMDL7xQntvDc3b2Q6CCVHuHoupwVGCnJu8QmW8Rs7oBtfxTJ8
sBIK8as+O2eCn2tQ6J8j40436z8LtkEQzjk5cR3/yG9yv6sbzoOwbqwPlO0Wzg1DEKal8IvLex+e
fu27jtsRb9QtzbKlYRm0bC5DXqdSP6KGp07TWt4ln2jhb4VDAqpaAn/+rpUZ0wot6DX1dC0bK96W
oZSrC24UQ0G2tghBCiEF9Wz7iSaBWWOFNhicKWMF17x41y9tDndM9i0rIFwg6G9OsuvdK/9x8YDM
jfjKcDA2R5SmBRC6odKICdOWqcQhqFT1z/0ONkIOpOZiFitSsTIpqUHUtX7u+TkCF/G2T3gNvfmc
QEe6Ohh01I8hZq+wJeIZjbzWDKYRwyPQ/AyszSC1qcgnKWzR8iNBycWd0+ZcZjsczgtJ3aTsYk8H
8EjEQzQXm99AfkaTEUwhSBl4TpiITZ1Ucel2sxeM/3WdBcJXccULnqby40VAQmeu2gmW0e63r2xf
k4qI+VAbvNtbnfXgR8YduKRbY/qv8gJd9OEx+1U16KycGikVxdxPtioVgz7twrJhqOt9ZMzg8jIu
1haWLVKa4lwl/qUiDJACsWPYDwMjxHf2dIwbuTOW5aH/xoo0fJqgf2xp1wzF9OFiT7/x05O7opdT
OoLVZhkgpKIKQ5f2mcFZW0FaGC0Bj+CdTLH8EjOeoSB/ajvC6tP8wfV7l9QlPloFUe06t6fdXyMs
vaZ1g0SFFslKzRHGTzVIHCycxeTpSoUt9DTBLvwrNKT7mHIYnMZuXh2GNlPMEK3RG/grHmmwB1JA
st4LitbsiPe2BFDKDPEs2+DBzqq62uM16hinaCYgEXwmxj6R924wiWSjYezZ+k3yqOG45ZJ3sO0c
k5olABcbe9AvF5aaLK3JLOLy7k73C35wr8DZRq+2t899zOrZCBdPTStfVd9Ejkm/VHNha/m8hAdO
wEUQp9+pypRIOQKUWstl3jGWlBjRdLpDRKBGf/O/J7ucPeL+AAYIYOLIVTFkZG6EsmjVcznKKyUA
LTh8U6+y5Sz7hRbXiUuXB/axOvT4LrTU29l9iVorM+QWukIcmJIOEEnQGT51WqO048tP7m00zVmj
uqw79bceDeEnEIsoEiWsAr+3ClTTUPMbzu9/q3k2zL852maFKthZ2mHUPoBuMWPO1kbcA0l8c8JU
hFm0sW+Admdyi7J/KhveelOPlrXMS1Xypcv4QFnuI+zaV940xtdjDKR9I8jB2nvKs6xsZCcFced/
5g4E0qXiEVXoXdunjGwjJWMWVOVps8v54cuIbS6OMzA+Pe5BQV0IZhyWjziO+kSHeSIjgvRpO9yz
lxmVl6Zn8KfnqsEJRd1oWThjEvNybsg6g3aLhwnaYT4PrSvpMIMbu38rK2+Sn7UkNzcnIIQnxnZC
8CwXB58iEIoc2dJpXUfbQ939PnJQJBDZ/Bo/QfbxtW5t18osw3Fm3CNOJA8sy7MLIWV3UJmy2/X8
+Eb2WGs+FS1kvo7NvJvEvVoL9DGtP1xl4NyLFSogsNyVEgwqwqaMXJ4KTelrR0Y3YWbkIPTm6c9j
XH9+sAbemCBulSB7u63fdjqWMfE86up2pmnvoSPYllZqcZGvUIWNi+i3UroWcofkGNjA3h5voa6V
KjnCB8G0nIhjtfK6RY0Qd6SmJMI1S/2dyWfOvbtMAq5Q7USr2bB5fitdO1BBmKhRZZoFVyvkyT3k
l1bgTHDwfehj9JUTVPOfdOwW6RHLDBudL7FB3cUnqEMFNQL8q8swobIWkTfFkWusAMz6fral7693
uyKjDO00W2gSkiqJguQlXFjDIW4MfTKAAHGyrY9Hq/o5jyqonq743K2ucMO3PmWWvVDkpMwwdfYJ
mIxwOPtRWgndoCgeH9P2aoAtuKnPC7m9Qq7yVWTMYa5Lsg2kS1a0rWJH1ur/RbL/Dva/xycg83FD
PV3HlOCFhwzKwPepht7kKdVa5HFF/yJu7B+QRLR3HM9OiEBKNYSjlhI5oep6JS6Xm78cRNaVs3zr
0El3Sea8sgH6YJee1AXp+B373m3ooD2DiuQsrILKBCWEpSdtKFZjH+fMtWbkU0O2sre/viT4ujhU
4ZKzdrYDk5OpjG7W2B9/e+ZADW0LUZdC2qY/+M/KZnIzCqEhLfBijuyDyZwmnQ+cFfxx/EvPD2mV
DldN/8IZa/Vigr4waqLPd7zg3BoUQHOymQFI361FjsHbDaGUS7OzHihtCj93gmKMpveFJYjgrwTD
Ohc9j/ECoQOVSc75PL/7C6Ub5CTUQbhBsKllNACIg+jghx9u3admOPQ2rAB5L89iEvHfme6n9N6J
UtmI7h39NQa4A9nSx5Hw1KX30GeevCkBwcQo1L5CF3am0aJtRb0zB+6lee+74TKIk+53cSgQAfVC
rqaifLLIuhEJc6TEliNlTmq9HesyeRX4B9Os3amdrdCeqd5p+zp5uCWgWfi4B5E4zttbKA50N7eZ
GVUNl0wFouNz1ZvkoPnMUWJgCFsKeR0qNXNv1i9fSIdTp3ex3oEMnmiYl4x88O+rqD2rNbdCNx+r
I2PConsf1B9v4/+RzprBgccUMJaQKtoQLCg20WG3Pht8z/WBy4xOGEkTqiJ6SHVe/E4Kxmq1EYHa
Wk3q9od8WKal/wUNFu3QnWanHpeRDKPjDMSp3L6rBoQeU/KSV7pBtPpS50C5oJ/Y7H6vs9U/myJr
08fsvwkyIRRZlCwg8SsQxAYxDCDuIRp49wj3g22pcQDN+XXJJ/oAkYOx5qCwHZ82QXtYKNEN7Cqb
HrjlHTYGF6Q/RwFsHh9NaStUncZgntHb10ItrItLLViCqZwD+cCI3SbJMVYgxvHhErHy0eyDuGR1
h3GYYlhwU2rG3BcT9YMXdewlapBY+Op1wclTc6hwSqiKkQM4tPWLPgnEM+YZgDZsQwg4rmrHii0T
KhaCoYKwuE6PmdRex9a0jJ/watqCi+mieozaekJTSv4gJXSxBf8HH55FnZwliFC0zlZl37RMXIqg
7UcXtR7cl80hUfHziHIi94Fc9sbpGHB9U4DNXnliB6x5wyarajijnjPbjqQGyv0988NXPMGlntdb
OVEruQqZfoNNQTZR+yQWaKqtQoEF+Ez98oHrmc2j8HpKS+XQrDk3VeoViuszDAv0nFDg1caBMkeS
LfBCAGZ5r/FtocgDkhTpOaYPfLF57+ZRXVCOfoWLqyhmF4LLOXUvlzbQjDfAVFn41qkjJbkV1mGR
J+7IYUOJ0Glv7Mo85dgIUxT/wT0vREcDwit6/owcsTb9hFbCfKQOqn7IJdCg6x7k8uMILzD4t7P7
1xWKLyyIRW/5nZHDo3EWN0DO1N05wICRWr8/NkzOfv6dotDrNSPE/YIL2kShHnu8PMojwSVh1EwF
+b9ml+ljSbPLdFf4BRIRGuuXLvXT+GvmT2eXXXEfu9Wkxvp8ZmIT45MRjDzJEHFrQReyIiYsabrj
ZFYnVFsVkF6osu8ERmOhO3jvKNYC7+CxPFDHHrbVmjSvc7edFwA+a6AOoCkmSzUDccv2Fjgvuy+9
EI+pppLCZyE5kHK9lkRDSSnGV8vrPqbKxDm+FGfawv3sDORh6vRtwhu/bFTaeZjP0bwzZVX7zTuP
Jnmnw+K1ZbzICamhj3qT0Z01GIVmTb2t0Vrt8VT2gr1JLS1pBhuLeMo04vQCC56T+PXKLhP0hDlF
aPS3wwQyVcm1VOYfm7WC75aj095U2+2DgU2IIlk1sIhEJv3AdSYkqX7Oj4+y8lDIDJqAWGeKJHFV
bC+Q+adsh9dil56Tbr8t6sdC6CJ4+byG2QBQ+druQtkWLg7iCZtnx9uWN6qLUIDZZkk2p9oC34lE
JXvGvxuxBHmfaj1Dps/LzL1i8bb4rnAVVp9gPb/TPeZwO/MCxhU2ZWhiUR5PZX95BzCtFZvabCdY
XUw63Ixa4pf3117IiX3Xm8ZjGJAf8tsHaWRR5uxAQnIF8CrW8OhLyf9ZA/Zsn0XeEWKH4Dwhes7t
OkNv+kYpI26MyuBwQMHYzWtzgKdcShcSaI/LzDgrrMyZgJBhr2TM4wyITUlU2KmTY2T6kN6l4puP
iy8ggbZ2uoRpIJDbz+3Hl/npi3VGO7UZKi6TXiJRQqeNXLn/KcQ6N8EvjCIBF1wug4zEAhaYwprw
cFqHEXQeGH9tpb1YAD2oY5ZIjlA7ex/QpjPTAqW545PLFKmprkCV1Yd9JzM+SeG9ceTUWCHEtWX7
ThQCy2DHIxbjr/IFPlx4k40dIvz4pQh/XoTMynU4GZpCB9TgIjaFFXy9BdU2b/cPez+FiXB/Zdmi
RsOH3h5YNew6hFILtc+IgWD4J5vxWu/NcB7Hrw+n7HIy5rB4DhXly+W2mY05F8g017l8PV3Ru1bV
NDawCE+vPOMpwAa0FNqGlwYB5OWxk9T+PrcfAOX80lb6ygfEP8j55YaF+oWifYAMu7fM3/bnN9Zw
cSQvzuJ+k3BNLnqT+XdsgUnipF4qmDed6wKYSRZWai2P5SODCD0VFxeKoqrNfPSGc2xvO40he0ZH
8nyF3STouxYGge9ODmRRvetQMYjvAr6y8HizO7xanb+Exg830hHtEgiAs6514SQp2X3epjyps6X4
CSK4oPv1qbVqp/hAaCJzil6tX+lA0XwXJqRC9Uc1o5sUbj1DUEQeis+80A20Tmo0keQ+W0ZMcjJ6
apfXAXtppBIWjZnAbRF6o6oh7M3FVCU1gE6aMFLdyKSYMMPoB/gng5DDmskTSy774AdqHlPgDmWq
NTC/YDKn4tKuYkuAecjIZpLsds6VExrpKMVbLqYrTivuWRiIPxGeJl/x+T4jkoR+K6LxE67ZEruo
xtsYrgBgVHdm98+oG8zBXKf6Hd7DYGuCeeLbDEgtGNzT6fYu8etb7DVSqhZBPIqli9kpFjzJtlRg
UCamjaKRyJgU7qtGpwWAy9TEj+6nSRMHnoP5NBVZzzmnI9+HkTyhLem49i1IGQKzVEPOhJrwDOMl
wx05WZF8MqnZ4SmJroY8dLZv6QsHafqcSpS69GgjhPJrUwan2Omx5c4b/L2J6tlCtDCW9JX/T09d
SRc4WKmdx1dkodzG4qax11jeRq72Ar/qjmDRlf6D3JwyGHMA5qfMrVr5CoI6Y5NmuX9duqgLzEiw
kon5AvBIo9Yuvj/MHoqzvRNf0rVrqLZCcVVJm7XZjcDw6aXDGa4TPSeXYCPzPap9GTfGXWgPRtng
g2+gXkJ2xYL1C5kpGrsPdF+00cHkpLEZU0OSckLh5x3Tto46YSMiH4p/5tBRTWOeaxWTkGFTTDqr
JEST/2i9SnFMp2vvpR7XifnRwJsElFQbHsYUu2uwm9VYej03P7vOh8lKG6nGQOp7NeNiQUMCp88D
zBgQ6JLz2HTPRzAHmTviB57lQ3ZNT42LK6K9g/Tag+5ceq6Uqs5hRRQG3fd9HUXBy1nb0pc7nxRT
20jBA14wE3OwS2a8w0/614IK/6lQMYdUljt2fZOEaB5AEOuylU35wHmlt2yB7V2ys0m0iWQ6wlQH
2bwo2FOzyfW64vp1nipIYDrZOthX8PQxpmqvJATxGu5I3Dd6D0lwQ3qBg2rUnvVbR9sf/AZVRhGJ
2kGypzWHsvxcsc4pj20qqYmxxlGJb25mm8rZ/59edjp88liQ31ThOuuqdPgdEJku4AmdMujqDoTD
lLqc6+b48GJBr9G2SB/zOWkI2e41nahAPByeWRMbjbiWrpt0tMmVo1yK3xO592H3cVjzQ+UijhYW
C1m3VeI2FFVWRYA/u1Ix7jO9cv0sLe8c38Ih9KAaY2Bc+/hwUeL0bkrYu3hiY1L7Id/YX/uWcHBd
QwtMZkMwMxWDeLKgsIQN/GMo4gH2rgplqhG27bw6cMpIKgjPZPOJaaqKLbd6VAtQTIGrDP2RBjEB
cMBv+HkKz1sfDq5u8c4eJTQMB9FwdLuQuij+uMFzYFctdFRTLOXGKCc4+tHLrjOM2TkDU8PbCUln
X3yx285s8KMk8UD3q5xOYZ9HCNjj2wPx4nN7t1WEzprZ21dqRyURPUplKI7Axdw1fDSfE8sHECwg
rrbHRCy1h9fd7EbA8BW6PsB1fXymDH87h4EvKhKm/tyy+7I6RcIT7ZuFiwXmtT8qvDUuiLv6ypk0
gnUGCAqQXKdHANhLrMsq+eczBZ/1BgQwKO/HsIlKVvbmct6UqFCh5RIaVG45g74gnbssTicVWoP8
bgl2UOAU/uaq52+QV0LW2BgsQJk0eufOeLi46O2Oc2eIkM04IaSL/jwpBXManun6koKltYBwYOtq
9NYhIv+ATrj/vgAiaIobdtLAleSPBneqUCYlM775J3KxwS0AiggwQvNnlNHx8FiBmS0rDq0wEWxs
pAb0C5cJzqz7BjqS3sX5S/icYfDw8jkEPFKxO/LtULiIwbZV7S2dnhrLZz5J+DICKxVEXhQQ3Znb
nEUjtPkOL33/Rbl8J3DLgdorqJ2ijrM2RKdIP3/Et/RIzXpz7/XSTueH12d+J1u4NyNjITdVAE/T
RDMOtdDZUD9p5/hOJUv5oxzIKvNe1pdr1jrCUCNYsn7ZDu0DPP9N8NWnmL2ofOWW/ONc3znjHjfY
fAwcUg9G/jY/qkXAjVeQMbkw49zob9euW1kM4+x4EdVUVS1y5oDUe/QTiRxZjIQiUoHPGX2Z9Rgj
qdF4pXUuWGE2fRCQCGQKuxJtYqZKCpI3OKOLvFyHxBdjiiUz6RDUbq/lJy3LQICa8eDtEtWcVyCp
b28wqZjL6szbNquGwCiR4ZABiQvwxGMXTBQg+6m2hEXMKorlH7HoP9QP3porpepAakmNCs0qYdfS
nkFPboi5HXp2dZtzm1Ey1/oPS9sWF1C9IJGBLzIB/Q+mMb+2DidDU20iWRxtyIlh96ZXtGpEwT+T
0ghl07mWd5sbBrtyN0Lg9Scz7L6atnhJSQAY/kccbcsVpgpby4HaGLFDP5Olw6uylEEQpE94Jf7o
/kzimplqdAKsmgB1SHdg0DSmiCR220HzxQkkEr4F56Wwc8BcXupZ+bt6oTmzdbwvEK2Kwioy/WpG
/uFMEINiakaE6suFT16lgV2+OXfXpJsppLDVE71BKicSD+SAJO52tTIQC+OmCq+3a2A8MhEk1xGD
ot3TBfeZxZOVq5A9WUyJ3LsiC49TNliC8EqrGCF3NrBKUQ0GhDGTYDh08xWYBnRChvg3HE82dKZ9
op2591U3iNJm/6qg8B4VQC9GfrFj9DrXwyBBJ2/+JPUoQneapcHTYdnIaoDIw1e2f37O4H/f/7hk
LkLv4hlaFdlsOJmh2UzOx/kE2xny4smfLFXYiyrambKI/eN5IUe+4MD4uNocJ3drrTkVhaEo5BqL
2OdAfzoSyL7LrqiV6rSpSh7cWtZ6wnjlbaoxw+nK1VrBCjQlW0kbmVepZCaD0lXPC0u5R4yBOeQi
+cmV+1SFXjgKzpda9X666QXtqXxuzwzkxYNZMJ9GSa1b7Ez6DfK7bmqISlgnK7zkWb6piOoK0ioF
lpViUvEIW72vAuDD1cM0qJ5yoKR4LhwUQvPzuRFPCyEcBWU86/BbjVkrklq4EFVQZXwUfhwK7DCi
SVyNfnJJY/rlYgolz4YIIA/W1VcAGDeiZAokQ18AFJW5yqn1f54vikzqEWsKBC42wJn8DxGoKGdP
NJV+zzPu4M90WG+6ffcBsobaFYmbtR4S5eYWypIuw8B3NoIKMwTdmusAGxflHgJhY70sMgeLU1LO
JYndFlZyuki/u+cJcIYwsgyah3LMZGMhg13+tQqUYt3+sO91Ptc07WDfB3thfuyS5bI6VJcTAIAf
Xlv7cb+afSJM8JY6MsONs/xu/YQxhIMpUiQnt6ul3aoGC/YgN60OOu0Jnf3YGoESHzB4kPP6DeAP
CHfsj23OyiCqF+r+EkEoyuj0jNf7d/PaIIC8JSXeQQOPn1/5iVT1Rd+kxSOMcR+28iKTaPRZmZjY
ijoBnmbClMZ3XT9OgbhvwMH4utzeG3ipXJ9HoLrpRMCs4Eak2kAHfWldBgjPwsAapmNikkgRM4NT
ndqvyIrLx1KLgfTxqKbF7l+6kaObu4ErBcUyPH9kRo5f54lhs0XV0aviylQUyZu9o7cbv5TDAuZt
ZSBL1UVEh4ZFUYmTL5KNSM2VfG/qzUexnrPNqFBMEB36RwnC0tVr4wL8dVUa5hYoNOb5BDtU0onz
9ckq9UZox1Ky8XZs5hUv3OtJ/cpt5U8x5Wjyke57Vs2B+StUbxBqb7ld0Dqnl85lNKMlFuabYX/2
pxNU+EKpW9aCzvXfai1YR65T4B52M6HJTY0Ty5hpaEM6p3P4YXOV4+VNLNg4dC//eHFdxSzoGHAG
b6XY0Ju8E5tVmtVR4NXqSr/JrAtpbjo0vX9sOVGAkkTgV92O2+ecoM3og/ASyDi8EkQwsJAIF3gH
IHpU58M7WrapJhyYVOCM+UTO2+nz2Q5Q2W7R/W2ncH4jGiHehdNDxpAAcdFcDqv5vSkbhYUd3aJR
OmkUJA7r68lRh32imvdiU6cUmW81sq0EMUHDfTrvzOH6+wKrDRo4m+m6xGSSUSJK2wRTFFul6g6c
9IZLCgbdAPNcCTouh/kUcP0Ot5+wZwm4p/lMFlhWC3w7e4+CReOLszBpkJA+qrYQbBBo5tb5i/42
7UP4TxnLjR/O0l5r1tnyMrg3nbJ5mi4RQIbCS22lFu4v1gukEJahTAuK7Gg+GUPPVbU66p/P5+WY
e/eOeW08lufcMYus4eqvu3MwAhUFGDBB0XDlckQMg161UtGZg0cRJb7T0R5Sb16axwmwNYOb0+UZ
DNqR5A1CwbUwWIae//S6DyKC3Gds6WkoptlXMJw0pgHeQOv9BrPYc7TtRn1Rt1oqL9WZAv3UBJYT
DQAAyxoBByZzXmSosL1I0LNvsScZjMo5IknZ8MFDb6+dBxj0V//j6awUbObnWh7fLBv+7Ds0lm8d
WtcARZXWu3Rssuj0stoSjCbSnwdXEMWQ3TZmizlrMOnjEhDk8gBVDogA4aTJCZ6YCULU1M9RvkAe
M04AaG8HuZxL7xK6K154w5e0NgXxOX520+6vO6Vd4QibYjKwT5PR6teRHoZL6rGCM3xogcaORryG
Vmywmh4eXbl1ip3n2gpsP7S5hZ5A1u297WCiHQ/KdbIdgNhCiiZ3M6+2+t3fCpR9tb4Wf/aa3WuZ
P1Q84fojed0Jh8AQpSmALYVhwTFT+1tjWWtLplSjRbTkI3R7OZsRJZSsYCTMZmMxhI/OkxLL85IL
EDXR1yAmRRt5/PPPBl/pD5MZGpQcks0tG5DSXYKAohXKFVLV2XC4DN9HymwN7rc/WOCwP16txyEM
em+RHzFDikqBquaLVIk4cvR0X7/wdUdJ4eWRUhsnRAatEBP0ZLxl5OV4PQ376LvzwXtx4Ul3HwyA
8/F6Vi6UHzew5OxIbfw8fM/t2jSr5Laj5cU9I3D9iYB+aSvhOx0xH4Rsofu7A6PJ3p51qpEf4E34
VxZGWnAahWYlvbkw8UMmO0atzp6gsrjjp6Ma8/X9SEzefaBSioCe50tRl7Vu0pYnRAa5WXQK52fy
QJDbe/si9xqXTaSvxsWvOlzRS+y1OENrVrZcXhlnCQdnmqKQbF14WkmA1bGRhUeFd3tBImtUBOMU
3S2GBqhBAC14jgMabFOPdU9P7X+3DCLNqG50NEkcgEaZF6oAchs02Knv3cJMAhzaCYn1kFgJWJz0
s4h+6WsJJMk2dbrYcZEi+0AP/0/rlhCO8B6X5/3HEGInICMi4cYiyM1wloFsL/OlVoL7J1MR6N9s
addB2RFfGWRbhIyUb5xRIgq1h/qee0y8EbmqYlty+zuSmEAZfDW5SzPdUFgYg2QBzd8FcQctgdPL
MpfoAwRUXpwgPx0vNZkYqGDhKniJaFLS0asq48x+TYI/FerW8s+F+MdDdTskGICUE4j7u9pYU+Xp
4JcrwWnrbcVLabdNiSYOCgNNXwdN2gic+WAJ5gLyJGDcKc7OBr620eHqzMre6Wgbz5kwlLx6irUQ
aqz75X86gwjm+hzCmTomFU5oL9OAyHW3xWuSF3/ZvpC0YdU99eXU9EpgZjWTAs8lNDR/aVOUJc9g
FiI/5TvRN/2FDK5f3aDaDXdB2laBT1YTSu5SzLsiG8wGkk+sl6/Z4j6JtwgSILTNAAkUL0t38cw3
HH1y4PsqUqg4Hh7VcU7/vRisLnfyml0AJGRLNgOdw3svZX/edBT4xNJybLWdyQrTuNMKyQKQ0cqm
yNVxJO87ke3lbmxbJOOP4WcvKUbWbNEGqpTbcH1+42EDocMTdEfTyTPI9Tq47dkqczCde0eklDJv
KApOR7x/zU607sUrx+qFikNH17nrMMVa95c8K4mzl84jjlAdyCfXacBMC97ZfBSVX1neNJsw4Gez
dK1XInHxZBJQsKQcb1X3FbzzvV1Ucwyqi2p2rcNhqtk8NHA6lxPBNCPpSlYczraqof9rSp/4oy8T
XQd/T0mF8PqUq/ZnikeVCNEUyfMc4oFZIwHgJgCFA3m2VHJucSu0Xa/xyINo47yECuAYT2mycyNm
XvhBzGMSTahyP5CorQefAA+ZyH5KUMDcI62Wdyv+qp6B3bHvfifQ94N05sUNg506rDQbAf20zIba
0p5HWoDKwh1D7Ntjw+yVljtFvfVMRnezcTObVprWxltezfDlUpuKn+uLXxJuKPFTVr8mmmsXefvp
5ODsFBC2BPP0BTkueZtm0LZsoWEY/KXa4heQ+PoanrY6pMcoSfXJuyLJUoLXaaLUVgNHtH2emKOZ
uCxxxSPQFbddlpuIGuqRbIxMzAtTRuKFoTouMUCw/BZtPqxB+rgJ4grFbHhm3YDjjhnu6lnQajDP
teBzK48GlD08cfq9Zitdox1RabEiUyvlcG08KfyruOrHwrY/Ps9jcuBypBr2tRsnfH+Yz7XavVR+
n9vR2ye9hcUdL/kci3AZO8h4ZXNGW7OVId1lFl9SvrawJkpa1sZQVi4yTh90SZW3QfSbO8/1k3ze
SpRVCwQ1oFytQaaAEjNn1YHcPG1MsSyl9hn66NeXmIBNHiFUAIhT8LAUckqO5xmMtPFzMsYmMNVz
3qAXoFZcQwwodwBYCV0GXQ2URzsoqLMiEh20ch45Qwjn6SuRTQbSdATHJzYT7k5VtJi9iIDql9xd
/f1MWxp4uCzcRxV9Q5Wl0XWfG3jcybLXx9rly3IFMqYgfWQm9H056uxu0jVq0BFcfvNgbDe4IsDH
T6rfUwxx7ZFh7T21/o84YP4rwWHsFVCk9tTF2I1lPY4ln1n71yUswB6Xo895pzsI+R0JnC+34HIL
JiRXI4dcb2woxHh67l3da5TGBYhPx3KbWWxfnbgMzvThMwRPLpJX+ojMuJrIeMgI1l9XiVvBn2pP
KCQ2HemPg6k/3W80OzxLNtN3ZidePv0lcqYmJU7EKwRYFpNITGmu4zTeFlWhMgYqAtO0PapmgDV0
teToYOzDZWjz34wn42u+Wm0j9cUoL9qZvN38baD0D9XEIeSS7qOj4FUYlHIzIvQLpCgGmzCtXCZy
q2vDmbZhUGfWQb0F16decvoz14oIPteWt5h19xYVVRXf5yntbuaBhZgZRMBqPZfIjBLAq3kWG+Os
XYsMYVn650BiH7votXeFivVXjWGbwCAaUTDi/RY454zK/368S1vYPopt14L9lLzaZxfyCnbyQ4Vu
RIt6b68cAN3owoOlU04jhF6lEewQhWUFefuVz90nMiBoSSWGFuaxY16vTJzHO6mrip3omEeiuRkJ
eWwftPe3NwYF5V5vyXKuflA16ODY7oVXLFRIvV9fE63JI4p77BwjAxtikdTOBGXuhk8EZoH1Roy2
TKuUnqaDlGL/YCjg4faOCRJSDEZtBTZXK3lweC0b1Bly7rVdsLtVlaTr/2lQO1A8tyLmoB+yA2wP
ph854e5BTKcUE/1fZrQhqR/dpqi1TefgTXPaCfkT2uBpCZCIEQxtjM9bbApS7Q5tRRI6QVzkjQ+n
B+X3pYlfWM+ODMXN8Fl4+zQtPk7qpZHRsYRSfL9jTQJZb+2efEns0ssovLvaZBj0qTMAFhRBhjMZ
rCArY/Qxgpfw4PZdO/HU9aifMjnQ2g2EEnsVJmdOZb4g9LxfCCcWWp/jsyKMLG7e2FbYqVIWPaef
+urqaMMr1cn14LGoCkD13PyRlHI1Bq9kZpN144JjWfxLznb1uEbWKaKAOqP00oMHLD3M2Sv6BIP5
6vs3rwkWRwU4JbBTlRvfoWAA/oh1RRhsqvNirXAPXYV1rpYMql+6yPtNyVq1dvbKk9HK6ibYh4fj
+QfoCw6qwGERGnKthvTh95a7xrosXAmpXWxFpit2KRVjGlNCiW3Xa2hoOTnJ/q5fxaCK6srVMXIr
CVicQR5jDYjZEQnBwmIxTMalMry+CO3b7EEqfezK5KOYjCETUxJNCTkUGBuWh1ojt66PhpNGp7WL
qGs0Sknjzlmeh+0uKKC27OaqKDc0oZP8wzM1h13HDSlL5taZB5yYcZMIvtMeLtPNzCN9QF37m3uM
S0oeoyVMOA/D23dh7J/gj3kDyYj4uGGLbT/ZGVE4bb/kufs0kto/RV7CnTPUmmymRBBswbWEcPdD
GNny7IDtEksr2JuBz4BnVixAvteNvQetuGEtzWWLwvfgWTvUJYsdNHooqrJkfy5+zlsL5gjz1cjt
y8KVWH9ygkgtxE/+uC14NsrBawJAaZ728QvzmmTcBhdvFC13kY3M67MZD+EWRFS914NZBaLOVyHm
H4cEGrKZF1qwCsCU7FxeU0R3I3wgEYcOA7zICIp6QrtwUfz3Q7AuLy4MM0GsTqHcUehyiHupzOrc
j03h01IrpSHh8GpiwJ0YQsAie1RNjI2Dsfov5YsSSmZFG1lYPk4LfS7u2V8/uXjiKEcK1RDrvY/s
ILxc1DzHlARZv1W/hGcNnwXwH/1D60Ic6oWyR1Omwb1arlFtVqqf798oz0hJQMI0l5NaYMdEnasO
m9MDKsUZDzgIzTlCsvpvsU517Ui64F3d4Byv1TMbV0Bo2+VRB282G6bIxlqP2G1x9NBZIiv8PLgL
dDeWxNIQuMT/fek0xIBhUQ67kXOlrE0f72FBe0JSCmVZr1wIhFHhg+hGAW3cLs0ZgKecwTHFfg4G
HZbJZ1IC56Q12+UqCfihcNjVxHFmiEu0pGVdeNcmqOsR/DEhr1D3K7HAJaMO+5u9aurbbX66Yrx1
horyR0OssBDbDCBrxFXLT+NNQX7nkzP447Q8q8tV5nGsTpkPuuAp33ArMMbnW3yPnMrCEGjWoPWt
XBzXOlWTj/SqNNmDM2kgGQl41hcdhJKDHDX3TynWWjuKMi4gpzcQbbD0NiLMtqOtPDTA09b3KIcv
nYSnDL/XunI8S073cCKxI8WSRnrcMtn4KvHGCI6JoFqyGQf+sJc/PCJavJtA3yiicPGcGo1XaHv1
NzXNdhmFeJDinBm7QU0+zOtK5yONbU2E/vrpxRD6gl7rQlovUfkmkO8JiUArO2IQimP1xap2E6zo
VCwpRlPvmhCqzo5TSSgXZxivMYytwHarQ8v6pcEgCvp+IDKGerkX8KeiPf/HnSRagLgEclHoW7ls
CA2o+A5JCVp0MCb1V5Tx+3KGSaW2xqdMFIcnfxcjxy2fDqmQtylCFkLQZJYvP13VGYLyzftoacuY
UpBAwOg5SXQtek+SCUJj8PWhysC/jhz1bCWb0LrE0ECtWgeySjwCDJa5H7SV4ojfs8B49+K4BRCW
c574WXItyW/vsrLogdat+ZlmxCmiYCisipFUjmi0fYXNRJhRkwdeOIvQHIw5U2jX0D1CIdjnFrXq
GVl62sIgLoO5H3yZgBjzKTBtKzPXRbP2HVTC04J98oJZPPuAHLLv/t9iZgg1SCZKPIJdYIFD096I
LfJlJOY4D6VinKZzTYbzFkH5ZfFo3INymun65jbLeodR7lDFxd6nqArku53D0im1Vod5JQd4NIM9
GLbj3WJAwxEgVwElLwRrLhG3SxLH2IUQ+8ThzIgMGK5ywoQIYjH40PoS3AkbZf1VR2kwmNucHyc8
zZ2aHoYU25dcx+uapDrhFM9I5p4iKDnyMq0hrgu4UtApmBnyl8j1PXgL+ktTDRYP+qRPEHNLvxNc
G7leMzQet1eQRTfCrJrVC7NnvVnp5PMEeVbODiOx5tuOCY9HMZBbRGO/ji2MXWCCu0Sy7izxijG9
Yo5NNLh0L9aUl6l5MX7o8Qai2gB1qv6mKjUb/UiSxLBNCRAsAX6Pbv79zfjJ1uBISSUdWFB7OhC3
ewbpLIxXcQj9noRPcaCNTKG3WJH29ew1dsmzJ7FbWaan404df1+gHLx+xj44mIjWDsHynL7qYVXY
S4VzfFTLWMWwDlsXwvcztEW7l5S+JSMLQsiI8TdUoH8coDThP2ZNq7HczZN6NNyGgT735Es9T7Wy
kuYs9fwl/TZysKpCA3otJSE64I8M9iPIYMI23pk/Yn52obqcuJqSIfshPU6AWp1/2pdlyGrIGx48
ncOCD0WrIBuR5kgHHVrzf0zedN4eHXy6OkNLdacDgoiVbaxVYJcM5+b2KGLWPyHfeHeFhmFv0+sB
N3DuGC3WY5iBzVeVMNQibJgNMixdjX8Bhce2P6KNe/yn8hSt1mdD+fDDp1sRMQASwXEu4dDUDosr
uKhHihUxbucyxOwpIG4PJin8ii4WOSNzhlVVg4lz7WnUGuJYbA0TloABD3+OChRkxfroXismtxrl
FV+Do2WdD+MRPHDO8u7h/TGoagzIT3syj+uf2mGIGI5m7kV19VNvnzdApRt0Aiw0mgSrFxun7gVc
vMOVjEao57I/fJVY6uW43PPmDWxng4ly5oxn/JNpFQ4jsFN5bOermu0NbR9XlFBY4Kv/bB32elJd
A+suu5bEgKh5ltENjpLj9udreVWnj5sfmVtsAKDmfx7si7HSkg8LcZ5hBvHOFbfep5Lhv7pdjAQu
z6fZKUFe+/m59R8OPqGg0xx/ISMKIHedFzZG52SO1zp4r00UVYX16XnBdZqucGEhvlbJsfnfSdQx
wXB/ddo9DVkdSvOKT4RoDYVz2uozz0iLFtqL7IT+Nnws/Mgs64wS6hb3L0ex2GqDdXgWUEWbnXsv
zz8gt++j6jp/1bFaM/UP9DXozW9wQoej1GrkcDac6V4jUWCondH9+J31C+5b+9d5xQqKyIsqy2Ea
615JNTVmDkMGmKMCrA1WiEL3sAtOp3xdtUMWjNl4jEOtQYyj9MChfHWtARYw1EfJwFelW0D6Vt8V
eSxV0ZC2y4ZdXWop38k2x3wV8pH7cz12tCI7v3WlktO1SSJCLjpeyWV5ewOwA1Tgp2oG4a+BxcUg
TrPnkfkLcebCaJjqZKO3J+TXStjgfbekDQZnljFwdGuN8Tpm+9Eo1m2MBxbUOkkjQh2E5J8bC83p
XbF29QXGemFnhyLK0xd9o30ODVdKD+lJ66K1Ow3sc21RNNwbsFojJdzaY1s43XQkd0oDchP8PbJT
4fv7PSc5qOfIR6wk1Osk/UMwwOJos7+JBoizrKycGpDyTrHcHVXGCZ/IyURJJnnzlSC9+ky61Rg1
x3kqpvo1RhL9P8SHDyJix00ge30Qsv7IbMC/QZpcL2WP0VX7MGHhkEE9N1XoKR313MRmLzeVakmN
/sCEugXdbEsDTpOt+l15FzxiajwMG34nsAubdQ77uzGAho9IYt5JxYR5lXmQ/CiqrxPPRgxHAh9x
bBzNlwcu+CFMA/A5G2DEuN2u7a7UdcthZZcnUFMTJyjfh9pPQRzoiyvpbG3iieC8KvibABmVLHh9
6Ti0rXA0VGRFK5ZUtdBQ1vOa/TR+cuQ2fAYx3L5/atP3MDbZOfBSdgmRZ1SPWOjeDAPoPZBua9Jb
zP5qliN9nb3m7elw8WxlI4hdv2oFwK0cOqCigp7Wh5vuM86dI8wGF0PRsjOBH/EsLtqJIzC0AOD1
WxuZ9q9ISQZrw0wStWOQM3RtFz5oI5ZrTHJU5j+YrKWLcPb3pXoolCN6BE7Pg9ZH25bW4SoNXeoE
K2jyG9Fs2jr+3vb0dncvT5U6uE7a9RAiheb/rZ40U9clH9Rrt8ElZWXCiXcadpRtRV0LxmtlP+kB
Ac7ig37ppw9R8+W1W1xzqpvaBS6g4vEITrT0BNk6Vro27PANiZhpOTLSlogVpwYn29tg8MFtazkn
o4ZTg+QIPvQN/3GGFHpI2GVIuCcXMaV79NG7LaTP/VHZKmkxMCd23TxtadN7NvNE41EPVbKilsbM
NEq44Pk6kKlvkMYB8XLVLtAHjR5WeRnG+3sGfnZkFEdyf3xv4/q7Nu2Swt6gJLju5d766SG+XUks
UiVsaCn7tTTH5omHZpYo3xvlqPVxBGr4Q/FSJkL1zYU3GraZDODO69/qwoQ1+Ze54JX4v2Bq3ZM+
6bn7Nk5Ble39voofg0hiD+lOhEA0qe5AeJiUzea77hVh/Snivm6b4MgoViULeNSKB4MJH6XOfe9U
/ZQm8HO8gLDQ5XePNTQ9CLPSzJ88uaxc6FWkowUGxZcsHmjPK3e1cc/6V9UT0HuW4qvsk8njkobQ
SdJlMOd+JCPa9cbQyj46rjBDXfDs/Z79LW6XAz57GWwHZBdkNQ9UARZXsNECMOGb1O/CwRPL18SM
01cZwYIhXyY5AxRzskT5uhdRp2wmKXT4hFd3b7I7oqLL2/eH/jKX1fMsTpXa4/l3qAIhcZw3zwh9
ygsV1l2rUqplFtuE+1AFenA+lNNpstn4tLqt/zq7GpePRw8oYJrMo3r5rD+SVm3YDxYgtwIBbYc3
uzMS3UXThgB+fr/QKgxrDtlYKDqUfV+SUIJpoCXi7+YWulhEDUH4WaPcJ6GRTlOzAqXfl2T4e41u
ZYjs2LQEHGRkpG8KY11dF2jJPfMeUAevCcuSz1U5XDlhswhGpHTYwdab4tXzY6zpWaRQV8sEktp7
fR9t9gOC6uiUX7TaoxeufEuzc2fmrIby02qXVXh6aYxB0y04xY454qJMbtEf9sb6Xt6RSqjyghTn
g8w29T/UzH/iWm2nDpx3XggiYLOYi0WW+pSajCAtPlgZKjhFo4alJACKG7HLaHOv/sqSa0CPjxqe
zceCRaZiGuTbcm5MwEcp1U8/TZzHATXq8tSNxZOa8yychsdyerVawXP2ZTbYQsXHZStsbNVyLgHb
Z6DMANTUV4NXlXplXYqUHBTag5onpSIcKjrpddpph05E9iHShY8deGolmonNYYb16JRzbiphvhSZ
SKDASXikPs2EiIy6fmpZM6wdTihp9slZRswZTonv3riXKLHHdLcvg2raG+tP2IfuWpakHfDshLWB
yQMxiFBAMGpqpNRG3OzK2gPnVxgAJfyer0/7+HDnMTQPUXj0H8tbDIcWuPCCiLIUvj4kZuxeltTW
PiMNYdPMcPSkeTwonZeTqSdCRsO4J0UtMPdVuEbS9IvVBTV+FbCDH57Xx/fnZ6olfHCSiHC5sEp6
+85QOYHdQkeCsRmowYa0E0dgJ6jm1sjARjFnH6uF2+bzzznn11434j2c3z7XQGnQbfTfRpzClQjS
+4R2Zy9v3z4x0bjMvT1ZWXGmhFQYqW0thoAokFDWV/ZYkKXJLIsBsRxvMRz9D5p8hrTQDv324yl1
eBwH8Ug4ort7GvAQcL0cJqIEdnYCxBV6aT5Ffcrzs+/kFGzNDWeMRd28uknA10F1IX4OZs3ZCOPk
+QFckn7QBk4VJ1gtXsJw+vQdBgUBNbtj/bZXHag5/sgzjn7eGq5HDCHIAUA7OpAA0AuTsNqcMp/d
fnwEwuWR0SKwDV2FElfsv2lWfPtwZAOU9BwTEoM/Mb1agwqJJY9Z/7cTgbtzU06EPZlmj5NYXbP6
VIPNZrpJ7GLNcAu9HA1mr036/trgPggKdCDm/hOaNg8c1VD4dB9hkdJT6RVt28zKqKL+4R9wXGLu
1ECUWF1Oz/Z2JW/FLKdD+CX5PcdVBE1sO/NeYSn0aowoH+uR2blefgcPu+VoozaK7OpyQ70Kon8U
6+qBDdtQqKaECo2980/Nevr5XnTIGrmWShbQqNFUWznL+ogCjZ/4vTGqL1ozAFKsSDf2YfXEP/e1
L8xU01THFYiZC4HJ5a5L4kKsrTd0zm3kbFSpxeLzJA8Jy955iZ8d3NaMGZYBfUhyve4BoyWmyivC
toY2jIwupP7yb62w6tW8FbL/HWA1cIxXUimtsZ7yXbU0LPuM5MW2WCzGnW8GJ2uHbDxXHiunm9Q5
M+0evBxu0hcpm9reVc1bAquS/c72ZkOqtX85tpJtTsQs8mxnJPtm08NcHsWwPkV0WOTjoRadf63H
q6cqOE2K9fcAY/lmkRREgiFamf+X5WLkY3+PyxxFBB9NweGyQZZ+ru+A6NqAnNqemYWmwtienzE+
4WJ+huBUhviPZ0V7M607dSfgPKt1VPrHfyovse4JQbzteTMASuYxY1qQM7cTmJBthYRdGQBFajoz
C7SEkSCI35v/8zNYNEn+Cm6zKQuuYNs9w0/bNdpe3kL1A2NBX02lvAeK4URhZsQsCYhGFcjnSJNo
j5wkm6TxIKEnX20/d0Ih9YLxwRPX9XJxWj0qyLj7zZYfWGbcOWWudxKjJf3Zg8mW8WoCP1gXfstv
fk6dzzkVTf/TB7s7rAkwC8m+KQjhjR14xFcSfiluhtfXkm4vm+M9c0R8wE0oM21yeakPi+8spQpI
CWYpVmLd59txcYPrzki04TUprEnvASpNeK6pHJgdCZLSuJgTwEPSPlIiednw/mm43sAh+LGQu0IW
b8z21pNeFEtuCRDQAMtlkjk/4iqBPGnkmx5AuIQq7nDJtgMjzIzTHzgNtj44ydGPK6PmyMmu2WY4
vR1dCCrlP4EeuPBXTA4SxFC2HtdPIsZNZvKcy98kS8jNqCNBV8eUqUYA75MvAanQjT0VwZnhw4mw
2sMbgO2eDeUCcKO8pwRDgR3vWgAlcDNDGIFN67o9GDg6gdT0vJbwErnQ11Rqjgde3E6QytyoXjU5
XpejpwVSWLwGzf4CNLhsO4lEcKeSnHNsKf79OZrVp0IQ0keiAyq0iNaW9B6ya7lTy3r0NrRj0pkf
+rsOItYMVwQ2c5dgirPJW9FL1r4Z2LPI20z+7t9xGh8dgB8X6a45v7bsalyMQTWPB3HCc+9tm9Nb
FJnsQsp8OynD7aUYkXeW+TRDthrePDQFY0DP542ADj3AG0KyVl4C2D6o7Uzm9vIT9pKEH5xbEGQI
+Uf4FvcAtJH7hHAqiFiIktYFU00Dvh3E1LMkW8mTba0wTCKpZH9OdZqc4c6ro0W/+NPLmrnMn6Io
qRivEDyP2aKsvenryESfyEA0L8XNnM/rcNjCWN804EmvdQ0fiCZweiPWTs3XCYRnj4qqCRerwcuj
PAeL5SSqjjYJ80l5QtM9ZddXUT2Uj3Yrb2jp/Od1CGg/ZmrUF4Q/i07m5JftAY4eL23S6jh0iVRF
B4Zil6by6JfOv5apCJnCit9m9HBQgIs4DSSAG1X/8+iv1WQsLxTniAHDYKKX0UAppPviHMdC/l0A
cJmc3fMjWZV7fbXAAAU+JcLF1C0b4yvWNU/Kc2mTJ3i9DP9wwtZWb0WrFV6gL0oHnTBmdeUs4RFP
iS/YMo5DB4RGR6+KAZb6/FiLrHf/UnSLo8Vto4AqMdwaWHj3H4Wdb5iU19gw0KtH8L5C1PnzjgZn
M6bHa4EoMFksc3gkgLHsGXwaGXpAYFay14Sqdhj0WpIVWc9/v5BbKXUL2VeOfWsoT3PIl52nZFUJ
D4cXa1A1e5K+wBq+Uibj3EFp6h0oZjD27eYOj1li1b2wU+XQu7jE8lnH6jSlZgYFk9486/Ed4iU0
x6RNAOCmBcx8yzxlY9Qr63oJ5BrMxqRw+JqUcLZ5BfBX5E+/4ngNKkI2eDaZQ4+kwZGFd7LT7tKY
2uFgdayfX8O4FnA7W7lrFNxApdbc2+Ys4j+BMD8CKnKuBB4fDtKpXeo4IH/QDpP7GmIIztF4hhsR
jTumdV0QucAIP0WMKYG5FV4znLTG6gouDIRtVjwgzlC9W1tWB/lBs4zmwZHw15me9cuQG3jlTiBj
evmLGmyhoFG/eUITg8SwHts4niAsfTTyT6+LDZx/RQp7p/9hE5bGQg7NTAJvyePX3UH0mII6y5N9
5JW2x90wzug8Ll88/QLhg//ceqUII8tsUhgMF3Sz5Wr0LRQgvCGNEY1tqXaQbUtw19bzo40VeFEt
dZVZixRA73clqKYZs6ztKwpqeos9c66d/pyN1mLYlf741h5NOP/CX7esLD+QdJXzd1HhOOpDAGnM
erMoMfLlCibL4F0hQDe7G7oDj4ka4igG4/z4PtbTbkICax5eyOl4pK7/AXj6oYk4CyK3ojLmjOJT
v0EceBkf0Cm3E7hDG1+ctrwarZVBasC1bJ8bK34dMyrEb7mNSQGSITDu3O1reOvPz7EZk1rlVcjd
t7ziyo4h+Lb7CTRQYlLDXGMrgGzKitDgYv7PgJJgCQ3rWvpt2aoVOwy9PuZBJLoWp1JCanJ3jRIL
7bXauVqPQzxwEbYr7UIrSd5U6aeEiRA+6geYVUCu4NT4dqrob9EoDvpIQT8SKCExk5jLu+eQcrX5
P8ohDkWblGbEcxW7sqxU7Blh7veYwNOMZkW4saBatRYAIjCbC5onLpnszPW01jgN1IUNp/OfYP0B
pPrFGbG0pLSa8HmUeoljEmlGSsn44o6XtoFRUi7GSwQGFZwDQgHDiS67FXeQRwahZd93+Js6/2zX
b1nVQ2N5FOTpPzImysC6a3EKUfWP8JVh80t5YNwQ1hyiHCsaOnApMMgXrKntSimx8ECDmYWNO0Ud
pfzZXTQFNQmy1bnSFaxMCSAaZbRoKl0+aHU/ouZXkn2oVyzgokB8f2zBFUxw8ZHY2dcdfj9XZcLh
sjHGroQi5nmOozFNQ8VDZsgTAK9ZITCghlKvZXMHLXaR15lsu/kIRs5Vy5DnY5W4Mu9NkBU8nYEc
klnsGAKVkyVgJrgSBuCB4kqyz6uJ170EY3ab3ELrJy3UbUXlB2gE402qCpXqDMj/4wlN6nJfXIys
MHeYGTavLlG57066nx6SSd9B21KOtJHaefUjZgToFk4pc6wEd6RnRhdRBlXTPZwcD/gdEqQMqoaK
onS2Or+OfAsA/t7QI56JoOAfRai2elun3aPU34R+PVUZ4qnPdEm3+Mq5pS24nH/0fwdaOjVGiDZL
r5vPdWwymQfZiInPDi0tcdDt85eOx3z4psKFCcsnuYCmD88rCSgnQcA5wApNjKL1PF6p7K/7u8UO
jH7YASjGw8r3AdmEjTXGFdC3gTOr4j60hR0EQDG1WL5/yYiOQOZePAZ7FufuyfTUotUxIiMmnSXO
F7nluLXJUiG9mApoWQMvTYDj8i0KfAlDBjoufg0lFGQFdiz3MgDFSZK1CuTt1dLWlQJpTFs1KmVN
zJpWylPSu+TED+xidGriKOzR1gS8GE9n7PDTsnE0ug5TCKU9j/nuIVmjhj7MsEOms9brlDdt6j/9
VtWHuGEaBXnMpY7vGVMahDLByk3WdeifvS6gs6bZGRSOPifgFs6hxv7AVcWiIcwJ3Bea5Ad8VVJp
0AI4Jre3VL8ndH362uHgGyicpK1I51TlqxASJ4pbnPUyV6dwO64VdUq5EdbrscIxHrIJnugf6IYV
nBMm/tdRTjcf12SF9FM8M9IINygkHXKeWD9hAx9Tb6hqgmfMyPwK6HdaD1V30mcsVSsC7D5J1Caa
nqWSedgC4rzCMy4viqCEtCK4HjxJEHQcztvQoEc5b4mfUAcUllkvQni4X7Q7ywJSxQitt6U0KCoG
v8m2XnG4I5pLM123tsrGP929K49x0nU46OHwkM5fhJsXZl8qMONoZbnno0UCb6xQE5/rVbYmkRFv
wlyA7SMaaSSYfivj4loYMa8VN7UyYPNlo38HSIxu4Th2GGsMZTUPhznszTy37Ch6JTZ1FwBbkFI8
N82K6WjboC6VRmB9jdgFCr6P88IB+J4TLvC+zn8GN+LzVhmBu3lCQ6jBp6aBEaWVpcFKF8DW4uTf
MJGrwbn7RdY8ly/r+PMVl0XrzvxLGFYHJjo8UkYOja09wFVlcai3GnAUmyJ9h1PbuQKq/xet9mv0
lInHrZSQTj7MZvKJvnrEeKESVs9i6XVCOnEhHZL7JSa8XUJe5wbO8c2Kh3qnuOcHsQ1xh064DLX+
6pRjJwItKHwaUHER1GOORrMi+bNoUmrINNZi93UX7sdqDWWUk2tEwffEKbsZCAfcVAoYKjTb2VmG
2wS2vKc8oTJNSm3lVvMM9D+cgTRvxafkNthWFFLYjHrI3r/qcvhDsGp5D5LDBjFmgF7LXBkOn+EZ
fIvGmEhrCrk7NjuL2YTKqcEFp1Hl4gtRQmFgs2npgPbQccqRCI8PvXS0Z6Rm99ypAj7sBw/0bM31
vjiWujnMF/C3TDkHv796WLT9wJa16M7ByJpUSs7iaOC2ZG7kYAdwVFmJi1Vi1yhHEYtYYwTZPhz2
kHUj1uBA8H4uhP3+gTYZvZuv5pdmh0d+9Ri1JSA5YzQp5FeSITnYkgRcqYk7AxG2+l1Dsx9+JD/o
mzse77OcYW1R3tYrm+DSP5swZXDS7lxg2W7vcXae+tElc+GAHeH9M2KGARwlocsO/ZD0MRiG3VEU
3qXVUOlUpRDbps1bh9GLZoMNDG3TOfKUNc3R1jfmdHbzTFr07RfQBPRir4HTK8Q5lcgThhYahkKV
wBruPpyHYkhIZEPCzWfrLh8dmJheTFIxh4QCtI7/NlJSx1qV0JfLG5iGsXicnT6gSNohyZOxwr1C
ehqcHD+aD/qmWwTCotSWYmbrotRVrneKIuhGEj/56EvhAwicxtTUwatnQxVJ0OBGGMtrqE3XA8Kq
fOMIcYjnY+9UTIVRLPBjKx7JOyICwYQanMdsBx7WmAtQrhE/ys8jDORDI9KhgqCPY8WACekLVllQ
vWsnSnKcw/h4e9NVgxvKHONvcF4LHrAaDUORYkw1acC95WwMzcCXDi4H73yVysahsRiCzkG1FiLc
E/pyBesdmWBO9Fb9EX4DQv1UdK7/MDskmlL6Wqz9kyBaRBgPIyn4SRjhb+twbw0LDX6d4AR3uX9u
xehamLfv7qoU2D4/HL44A6IjCp82ZjhFCsDjlX+tA4EZQN2wnJSuf4sr+I43btCwzd3U82cvKLjy
ZCEzpZZpQpo2RUXExi5MeKUwxnKc3a3KnUGKE/KvFnpuBU5RNvaBkW7ukUa7HNH3J0Sp931Zv31o
I7pa+CpdQuxuyUdAFsWx45+JMylbgnc8XkyG+O2sbk4POMvDDV9HqaQ6rA9t/fat/HwOHa4ELxsd
xHC+RuZh8nFab8+o+1wLMsSYkw9i0Coyg0f+3Ekzybu+phjuNDU5ybAtBYXFToURaaSk9kCGOk76
i4OufUi8jR+mu8M/rbiWY8am2JlGS3Gsm2Vn79pptszmsxeviV6zH6r9ec/Je3VBlW/ZiMRX43qX
Vs4Yo1+L4Tz3VwxU8wRBL5WcUBfZAK1ylrZpFTRSF/zJHkG/STQEfYmJZcaNHuT4/ExhZ4EBBjSZ
TY+zjqvJVYSt8KcLNFUIwgND/x9Ujp/9Gzyn5bVq3OyKNigHXg5uf2xyF3GuNLoUqguyNeYV8t2v
JD84D1zKmnMKlkJhT5CvbK+U0hw8tfTQegXv9mG4LDjvxJb3+EUOte6NAf9HORgS4lzFBwx0O0Zr
Ya7oxQG6yqDZQlbgdtogDfcuyDX2zGGzdtKxim0TOFzfL6M+8MZCqk7XyCeJ5+M0Uv26WXoQISSm
ne6J9tSA0KukOUn77UMl+KMW8KuV7H8SzDqcAafAAHhUy5GYeCS9jhkwjy7OMb954e5AzOfSasTO
0nM9ZFOszFF0b3xjlIJFkyKblePHTG4PPeje3rfTEzoxTZGHXcaLzPpkFLYpxK4RqZu3FHhScuNN
PtHVfOu7m0bQMBLKiSIOCGHYYl4v0MihLvs0usHJV3EDFquGk3ezpLEzqlB0/koPrquD92aO96lE
2402as+Q7uR7eukdC9MRtzijYDvZsGqM5i3pyEbJFx0w78w5hkxuk5cnYnPXKPKX5oc14tlPkrzQ
QcZ9oJmrPzvu88y25VWQB4PKcliJ8Fmwl6D7a9IRcxtYJqHxhUSe5FJ3sKRCKE8th7WuDuXZPuw2
Lyk4hKRxKZ0yQiasFUe9pwJrwZ3vA+/nwLFAiFmO5uD8qw2N8JgbCzP7PvPQ3Ck+TUjthCzYeR+h
h02R/dELvaCVLC1LLaTyEp732mI2lrh7TV2W/rqIPS9lx9r7yFu9uCX97P6YNNW9Xfzo7ogD5hXq
OjKcK553SofY9WfvjOXlylLMZMlcFiNBlGCGefBzUOsA4kZH/+eo5UZR58o5p8/OB6UzLZT4XeHy
9vieOrDoIShXjSkCsjLVEEIUsl4imlAp9XtRHHafiDavbvE0mBEL7qa2Gzykf4njmWRI1SEZfXFK
PLZ3RZcq8wXeixz0oAs4O+YfXT6rkbPQhCGpu+ljFV0lKzxLq7FdG8o2SA4jKuq2C8ubusAwNXNI
KOXGL9LUrifR4mdSbEBLA42s2tW/c2xHTev/kFEsG2Tmz1syDabiazFDeHUTBAhmk3vYbLTuJucU
RpDL7RRvvW6P7rNKpT46Essvl+dJR3QRc5Q9bVB8g4yqL7A1TgeghShXTVHJ7yNtiUgRRBELq4EE
4rc8sJ72npLuVyv2f+GQw65vK7TMKqJZaY8adH8KJd8rZ5vGxjRqYmXsrL4SiK/Zfgrt7Sh7WTGz
bJvWaBSpMRRDAwzlHpTgU9kyL1lOa6z9UcCEOgmBkEBUEtw0xAI1wYL9o9ujrJfCRyzXiqAQYgKh
ijw4A525GP2s2yjPdKqI2djkeFm/Eo/SZH6idghBD5gIaxu+4gvEz1i56BoQoZpvsPVmQ6JnHW1D
MKpqqQOuxUJy2r3VLIQ/K4HJ3HHqJ4a7CzxKb9ImUvZW5rWx20Bs6VrLNIz1nlK5bU10e0tQrTe2
q6RXu3+z3QYq2Rivx1ytyvEflbNVz9QqVTh8qvGF5DcFLoMeaXpaQ9s8iQ/AwgJqKhKQrfNfNBsP
Jyp9l5QQwPkBW1BQYqDShoZC/GUA72uuc4pX4DnLoIk+IFWF1twnhokLxegorzbUzmwVPmepkQni
iNNPGruNhMvvgZht/ye4I4Zyl6S29n65nKnTBBv0f0eTHOJqgsyDt8rCuQJ4ijavNTRHdgXLFJi7
C4X2pxA7oKruiDd06LS353Z66DpHm5GujDqf/7B2mEpRo7fV+x4x3UZEXJgiqPgyF7IkwyZeRNhc
gfAP/+VQAkItTfSVpR9f2FkeymSa8YBpY6Hl212VKSRb3BpmTTaWISOSdQOJKv202lPm6+vGEHOH
/dcHYEuv3I4ihffXqfyshKLGiZxPdof3yAFqvkbPKYVKp1fbTDcfM/wj51prKUvItW5qSXdH/Vr5
mO+1k3OHzxclcjXhEROOFGpjjvak1Dp1aNIq79vdar346kFGnVlgLXO2YxG2nVrJhOvwiZnhmvf5
wg5TB0AQ2s8jfR5TL8Pmd5+SnyQKkE1gwsvSdjcArQe+SjwIi4vcCJd26R46M+3nxxsAaj+qiT1e
bLhotBF7lD5wp4bbKBGWOcU/lxno2p8lGHYghssmVtP2CsnPw6O28W5ok5tNsj3SFZMEJANQm8EJ
GQS2qjnv0SPWE1/0JG+ORKFjm3S5fLRbNYZPQa2/g04+ubb1klQT8sHZcimNMPeE78yFxFPIBYnj
0aMxl2aW9XH2BCk9538d4Fuah5VilCD8uHZgYxbg79mwPyTWcuDQP5/HMVHQHx/DJMjEl4sK96MH
vl2uwI0ghj1StFPhVEjvzDvZLehoHgH+WWakK+86JIGhga27iz59mNRQY2ZaDzkHx/ixKVOu/iyG
zwBYnf8KwbIhfJoCEU9u7frHLapjbmdHE8D+lwT1a1p7N1lB17Mo+p4WqozUylDm8Ok5Sv1WE7Ce
7lls+akaJCUNL5CTri5HwMmN3C+K1XKQH1N727sasG9vdxjrY/nCOXNr0qOEZU5TZxmmzS2dteZo
XygVqYx3P5S3Yn5GaSjXtOQeJk1ifQ+QcmhyNvslw88KkS4HfESbLjNFLOBsFgtuN5yBmc4cKuJL
yNBQkvbAZ+cL75j5ouIevZWU/vbhO/r4tA9sna0wdqRgaaSWc7ci1rV6aWH9xlRekA9qITmt0ZTC
LY5wAYFqT8Kt6leCoj5qrIWIxyp0uL/odlhizh2sJqTevuV+UXS8V2sdY6bxVQ2pjGos6nLm7JPx
biXXRsNHdCclORKQH9KqkCKvv2S9o6jtmisS5kyEWqpVROiMXGIRLG5Gj5Ka8OYtWb8eijExl3vI
m31fWweWQXba8+RCio1F+zSBefdXIuW8Cgr5Se2sdk0w2Aye+6XhT18YrnYSKceWmpEf2SUkV9A9
Q39st3fiqLovezczyTBfF/JUD81qxvDHtgBdLZcvkBVINB1PbUP6sGnijbDOnK599rlvM6w4MtOY
7CigHxwONdt71hvtbEXCA7vpeKKGjoFzMMDy4GIOZ3vL7JBA92gce20gNIjNeYP0XorVjENZy6/x
v6GKXBHuZKmaTGQj0BXDYwqQT4d87VHhZXivP50654sTOo1n+zseH7cUsykQwS//p9SNtsz1jVEr
F4HVb+OuxdrszPEgOKBZQnh34jETVDbejPM0Ta+ih0BM27cuiNbTWIdJHWXX1lghIE0Wv7HhPPmL
eTkD0oBrzkJ4I5KawyNffx0hi/dJ7TPQrSMPPu3am/2klxqpni3Lw8a12JKCvlBWjufKN8DBdYHm
ReW5l1ZknZ+ooOfMKjKeSEZ+WGm+dpXzuBZ4wNnvOrduAB5f4IasvGq45fCKjfVpnRMTUl6GvX1Q
Np4C6lK2TmPRayuI1BGjYmlcsxewZ5vfGzrjSJJq1AvsKdT2r+pijj1CN876ovhf/avOn3l0xIy8
nB9AnNOSTufnA4on5e9Q4AEd8duvBADPFxu4FC2cIgLKwLdATGO6uNxOTlSEiFo23N8GvEki97WK
QD5DV+tbI85GPZMdQOegHl61Lyj+9DOb3XjGaXaYiyV0orBAKyAX+nfxSqWEJ2e52DIxtuCRZNJ7
B2/i0ZdC07t7fKF+4OBqLd6I7gyvJj8SP85882lk+2FRxAE8bMm4O7f7Lx0MXNaFPAPta0uNTQ6T
JiwrumVGXUJSoaT5rr2VUu2/ThGjmLfsES9hWIVIovZedAoh5Wr30XC1+tbC7TRGDohjT4+s9M0I
oiQWE3WFFc0UH+aNAnp4zixqPcFXipjTEBlmPZ7YW05lVIxoGoBTvG7m53KybGctULIomJkhnvOJ
cB+feLh+DndCvriYhmc1GI7NlHGlo7oujBoFLnaFdhldgcU45Q0wHbJc691qrEdsfxWp9lv8pkCE
OuFIWYtBkEK6XoRHxvxNjXL9eeJLz6v3RjL/SM6jKQZCQXbu33QR9wjvVn25S2G5DtSMagFTToDp
Gdx1espCxRqn+m5qF5+tBrkmsKBirj1XxIntB3a83TTk9SVIKiJ+3demAMtb0XLKpZMClmOztuFB
G+HAYApo4ywpcOe/Z1A/luFyNWEfS9Wlu41ogWvlEIOMLhstkklxqdh5bISaNyAUSWruAIwGlYYk
pzNb8vcA98gL74SIL9EUj47jMowYFJdrvonQT+Rdh3/vi284BoS4hkuOgJ20OkjZNUNJ7a4XN1Up
nJjW4AnEtZCx4INKnhDj1oyoJwzpfZxUfy+k/+wEVgS45oKjw12vPxjfjxsMXq+33gGVEicjARFx
zSy/JXPtinN88e0M4hEgn3ikDa1SDlENIKzg0IqgPaPe6HRq3nnRj1A3Cv73RJAhOYG7P/NYU78t
3yReQkkByTNqm/Q24BwfCOsYw8KuoaYhB/FtuwXrFl6K0F+yX9SiMUPhMrs+Z7eqpT9OI/iRPY5D
4iWAeMImsXfPV1F2hxEC0AJ4CsL5BtdNpF5EjjiNH+to+6skmlxIYs2U5eA3ayXVEYF/TonBh6NA
/s7q+y1dlTwXnAoSOOxk8r/UVmaF1KjJ6fmTG43fOw9kjJJhq3VCujHGQcnIOWGPU9lVScKawLSj
pwjfHUleMLMvcSuad6fo8McJNFeVIZPAj9B3XObXiUqOoSVdCHcRogYg6xXS/hIWbJJpynRtD10m
uXMp4JrljcadWeEQ7B4ZHEDxJruQGMqOFpduVFDWn3qpgm2LrxNzuGPt4O3AAbGQPfAVCBJ6y8qr
jWRD5QLbWzBLwsrkAl+gfb7xo6G67LFFuOlTY6LZ7tJA8+AEuKin3St8aQwfsRuH1dITnXN7BZh7
d9beVPIwSeOz3mUtyXtlwSWNGBNgIhMlIso5q2J4wj+jS0zD3HKkjqUALj8RNb6+TlVL37PyFgwv
/f+OTWbXBWq0zcOx8sjn0W8aGqYUdL/B8lMRebEYC8RXPjSRY5coOtZqLSxWDtiwci4w7a/k6TVU
qKhLxSh3Zt+RidA8Nlaxe8Ex7nElkZg7uy0XMNlBdolT/8z6wisly3oH9TA38wVDA2wKi9oxmJQc
bYOyX1KZi0XYYJaGDD609Ew7lhF4eJgGBgwsVP/MGS3jJ7BEtd4rG2gyYtOb/qsr5jrRLvHU0bNy
t0FMgsR/8Y9D2/c0ojxrlG5bRFeOuAkeDN9zB8TIV9Sd1+cGz3inqmnrfQUbrhZptcmql2fRSWFY
5y6yR8ewHZdbehVEklkXkDP4IjvfXZTcFPJyAdOIpL/7yYKq5v3Jo6do38qa2u6Sctl97Bh0eSnW
4aHy4lF+K0+06TL30Ufvc6gH+Q8bef8AknOdosS1P/b3ZKKkAuGBepaYO0mmobjQhdE15cBTGf4J
IOsBZZvho13Ena3Cwq/Hv2YvIqOMDyBGgknzezcd06eCAIQzDrZ4uln5oHG/kSDQZHWBwkan5cw7
frzpWCeCklxByjfs+YpAg95wXZ1lolg2UNdESOaS+sqyPa75negStvaIfbykgGS91+A2j4oZIELm
yUOWEK65xvRxi/KMLqLSO04hUwcLAhWUTkGPUtmqbrPBswM8j9nPC0vWqU9cBPVL6pdGj8LoqHMo
5autsBK6DeAvd6sq603WrTez+T3whxc/m+xUUq+nocLuoVxtJ3iI9GrJBbK+hPZwGcrJCPbwfB7I
sVskMZaOiVOe6dCIyUxj98Mpha5nFn8aF9sSUiLfcaS3eMg1o2Y2jhVi1ejzwVMX8wFIJcuCvWyZ
euwJOmu3URGQwJ3mnQezZrl2wfSyKgbsM1AUlJX+QUxyPNcIt0sO6IFzampi3ZEbjOsGHcRxZiPr
3I2ZsAhti28p3JbpZXvv4AhJDCdP10lKBYgbwfKDXX/WoAf9+0msP6IRbtcSMbf6jNai9k2li2x5
9Efls0AO0dCOjVOpq0bF6fv7eXy9lMKO4OUW6azgBunlud8itXu2c+iMivdVy/9zKfeMQ5EFijiz
+W5xD7p/45VsQJjkLtIwoeBcZPITcVaQPGakzqiC0d84gEUq5Wf9t99JCfKo/MLg6JLzRmAzLotX
D9qod/GolK0Vm2ycWG76/+4oPL28CunGTd7DBD8BuUQe8qnwjNarxheJYnpIQdioGZesZ6RLCQLl
Y6de9gJthMdqbWqX95LfRhL8+nIJNWksMnp6nUAEhijBXT9q9sRnj9nhFT7ecvg/+tloIWeMJ0Lb
SrALmEuiMpDo3u7ZEXVCoYuqyP8KLnx/H99viBI82VluEoqn+Wstqtsz14gwkxPZ19xvvkuxzNdI
3XBsnrI6MrULavfWf//mpfceJmg5QgGpYUG/SjjDq3UuFGvv59M03Qitut1txQjpS4nSjq62gVxO
TMF7+00OFsfUFjVKyQlda6dAH31Y429bihqN4MNH89fNxMJkek3MjQHFFB2FUMhv3uXi8RYWPmja
UQ3hiYBuhJnIzeyPHqdFCYkiOljkN45sS7n6fUw8igWt7Ys4lIvTfKA/kaKm3g//C6VdvyFLqtRh
EphZJ93t9ItpsHxYvs3PKfbi7X1jDDUlPLHhnJzRHxaqomDiL4e2MjslVHrCAf4HW8dkczWVszCh
JcJfJOPNDY0haJczso0qTw/6Rla2IubhbTWCiDu+jQs1sjWljaqSkBjlOYVIouX3HgcOevozKTOr
7riu2JON9BAjiAN1trln1YlynRbeek+YsHZ3rsAITBeMJf8qsH0UVAkvKTkQW9mC64PxAepeKwyd
UzdanDu/3wud31ECbWw+34yVl9kEBpts847Brx1duL68+652H1id333CzAWfF3mHCnk9NvRGX/+Y
4urxvoxXK7jeQdnEgM9sxXf31iK96hpT5tuwyRNJ6+aJvMMJbWCMEDF4/Z6RfS1tgUnLnHeGtphN
SFGMSi6RnVeXvHPXyHSjngOm3OAe+ZYbsZHEoBoei5qd7fp/MWdTRSFXtVFFWhWZcQzQU5AGPx2q
GecESiPBi3AHGAnuHYZNpy5bqQKJ5TcJf6QItyatt2vXlyBacbMiGMkUgEo0SawwG5koSg6nOxv6
B3U7BHM2Xk3FZ94YPcjgtax6kLuwOCVKMGonpXj5pOLBgEwWmTRETZKB0TEfTbnYQQRH9kFJbUGf
ENbtQZcvnwAbiAq1sr17CG7V1fsQ0/hrxCYNKbJfixaCSGkM/TuHs4Goexh8SZ2c6/Od+xq/JbLz
iTPXGDaPxskkDxFhyg5AcChAshI1Ws/LuRZA+/j3cnUgtPRwr4DCst743EfP/cLE8p0JPfGu5uGq
0JxNMu4Kjmh/+GGhdAtljkVXqB4u00jO/rL/897yzQA4YZrqPxFkr/01ufCA6GeeIby3rH227dDa
CCkDLuJNmUM3+e9pFY2if5hRcc+S1zXW+xkmZdtlVFmSDQ2/trOfdGOF8mAy/lGZ3NnGg0twFcRN
RiB05JT6Puad7mMesMusO5znPB1emW9q9eevY0BNnocgsEtVBkX/t0u4nW05IJxe8R/s4R2/lhft
9yyYyrJTNkfyHUDbk8zH9AT5t4vlcbUHwsOFmHMY9eFWnA3ndUB7qs13Vg4aK+ohs6xocPPv8xbS
mxqbKMY7i3VWmV8gvESxSpH6n/qEMmDEbiDyql+qPtEktzIW1GA+iMyBrMu/dwEQPN0nLSAgUIJ+
Pf7lhCiCjoGg/xnMwGDMMdfhMRt01kDYYMbQVGRfFfPU2dhtiVgUiH2nI22CjpsTpWNasQyLi928
Hb6Ge8uViMLaCJGUlkeg4gsUmIthNH+aI2PeDeO4Q1uGigJaWUPewGm70Zg5a0/3b66qDuo+/8CH
O4qS4SzxWDREFCNZhe8MCOFaPO+kwHekXsACirDZ6bJc84TpRTJI+5tnurZVeds4e+T8d0UGztI5
Sf+OS+ctzC9ojBfa2USJ/MZMQ9PI+JBS+ofiwPAgk9uyY+M9Sx9FOpfjFYoytq+FFT6PlVulzbfY
9YiN2kdElE1/CI1J0MmsYPpb2xMmbdqId3qjN8eLkHXhxd4fHkJssXTW1Qqv4fn58YpxW0FTn7nX
Jh43l5qmlKWuIwjj2JU/dD6X/Lkf++PRQB/WZn+K3hqptza/F7bXMRCIwli3Rxik92NKq+9NMdI5
pfFGoi7PFO3xQRGqRlcqTMyEc5YhtYFsbHVG9DUAEkvWaMa53/bt91WOaQLhEtcLSsXrwk2f02Hj
h877B6VvulWoyOOh40b+tj6VZXv8kBOKI2iX7fajCZ8Qg33FI2OlHjF3qlz44m+k80TeJkgraq6G
VxLJuk6/HOkgV4j65tZHmHFnoO03uafXcTkWO87it30x5/Bt/mfISbcmsT7/7KNLEcVpm6XBaAZz
kksjl4WfDZyIaISZJAEPpua+FemovEa6DnZDuIccitR4lcT2zduuTFRYLJT4qAwYYH7MITMh7rFm
FF7+CXjHYtobV+NSWFVSj6qWWW2MjYOnsL5qYr3yAhuNHavYAzGV2tjlfy3y8ndUEsOircNa4USq
uhi9qP9+ue+GK8nMjSRIkjO/mUoA34W0pmRD3KWs54GuLogjhSeAurCQqoq88oGOdn9I5uynmH2t
AEMpDtfIIGUVSqAfkzlqsKsVZ3/kjegZegwRmGhV8FV7Sd5rdkWejYUQjp/kHNBUTDNyZj5q/wvb
j+MxCi/xV4xDhON2UfkQdLw6ctNJbmoPVRmsCuU9+3XFt60Lz2PFYm5wZGGuFUFKjPIpRIGJc4dG
QDC8muNE9osXRGNEMziWtMy77mX0YZDqAu4BMZMSHFqRQ6kaSBUh37/ccGQJheZOffF+U+ssEx/c
if3dYjMFcS68A6kAAGkP91Xb6Xc7qd15YEwUQbGXigrOUTWs4DB80uFUjJuFLftvLH2sMMQDYiN4
lQlDpJO+9B1NVw4AcRLItnbvEDZpOMehSSG/dDqWCUSkHO0qJmRndzYA2siuezATHDTvvsZQcXL3
gryHMDPmBQD8y3p8B4GLcqU7lZLNlsaIaimW93xUq2GvoV9UssgCevE4o2MyRRh0vFw+Kd8gO1Z7
MrA995PTqIPCnHh/ypk0XPWgxUkBRd3r3z9EH/KF4PJrZCZO51m+XhhbS1bFfIA47AutKKFhdro2
zhgDcoWFYo8rK9tyqUfXHcog2s6dlD5MN5gIcHJ2d1T2cjYQusAC5Bi1ZjcIhRUcAB8tBhlGZ7++
oBK8NO4BDAQSx1SsU9aDknip85PEf8obF0/c7zqQlO9pUwlVQZn4/jmhSerlzIKm0/uNaQtbSoDH
Ma+tC5zLX2lgz4SJBEl/ahkqZyu1a9IakPbPC6UZfiZQ3k76BYI2cDt+idmja8mt2uJ2GySUhUhq
YEmQl9BdiC2QhDUficI4efpW4W4G9fpdj9FYj2DBWNRjH6Xo0XPQbi0cyzF4dT2ii9vZlgBixycQ
olH2YiJ/67oz6nr/sEfsptXM+wiC4d10dXbmorJTuYdo3WzDp0R4t1Qf/vqgLI2q2eK4qK9Rh69L
e/zY6paEKzCR/uvu4zK/qcF2obBT6UMNk6YGlP8nT56VPEsjdBQuHF9I2qJOSNLguE6BGWHzcK+I
9ZQSKfAIoz2wRaJ2hfVDf0Bp18H79OZswIRkr6mlqXnA7KUvkHqxXUGwdnO28H1+ADy1nqcPojHG
TFoHfubkMsI5HMx7g72S1Rl5CA7kdSSyv5ybPe7Tw9WSXCqGcVIuN8stoTuqNaAFEdd/0J3AgbQO
t+mO7oh6UytF0JIp7t58LPnoSyMpqJs1RLfSOgJ08WnLeGnYW5BQFKXDFqr5I+fNHT1hpZUntGEz
m9BjObGFTpBX9CcyY+7otRZFi1dCbm8c5dlXxNY2otCVraX+UYosbAuSh1liTIWS94GCBIjWbRul
sSF5rAzVqhrUyyHcfD781Ql7jTleltjHuM5VTtXs7EzX0Uy5tsHEZbxAVnrQRKzAFFvJ+sc6HKN4
qvQ7BLFR9CNLkZrbr7g1+c+rZoQctY4v0NagXFybz1NPn8NIpOgpzRauOpE/q4YEbbYj1B/87v5S
4YL/HCUrO5O8YMnH2VZIJTWbxBgjZpBNghHYOiqQ+2HTL4r1Yc/3OjyuVO3e9A/BMQTua2Uz40jb
CWzdkXhN6kFiXlNgPpqWUIuPn6Xvtk01V0OFZg1Bj0PYNAYz8fjMhT0AFcM6pYpdM0eHOgnvwUGe
gkwdeQbNtqVPeTBC0zn/+bJ6Duq0JgumFe19cxrqhN67WMW836mI/0yD2oFtuos8tE5T5b3wP0BE
DwxVBtriXHsYY1jB46tNxPUZ41/b11K8HU1Idcchsbur21rJ6hbE4+fAapqwsZKG0kEV5FU0tVpw
8+shpuPeCmbyrrJYFS7gl345D72Jaree9uOxgS4CiDJy6iGkA3KnOWpnlPU3na7XEB0wC62N4/6Z
5Og/RNVUHSzP9F8qEfirijzj75AONYtnBIogBVWA2zmqhK2PXRZ0k7GuyhNMjQyL6RGn5hknoT1i
EEhwLNFk7cwQQXfMqhLkrtiP6E+hxBe4wiBW4BLpmetwBteWiEupRuOwNfZ0g3J2hqaVHuUoq+G3
hOVB1sIvFrErTnYszTSxae/gI8H/15s93z2ixpJ+WzDo/9Uy9TQCHWioyRlM9Js/Mfl4682ZNKtM
IvSbiG0es+eF3BAkxKuV3KXRDv/JTYdy1bd4VkJ+kdXJ49ikfWfd9+CFikIXo+/5pNlOYbSEDoXv
K3CCbJH1XICZwRT4yG32oTX3UF651vPSszb9T0Xjz9Nf8pSavjm+9e3mVr7nK4oI9SRdL1coMjHS
zbs5xFyjSfpAzeDmiv38P8ILqbQ5VKy9uSzkzPVFQ5Z2//McKfJ+bWOYf0QHze7MuaSYFr9BXVdM
1U7URj7YZzNtaWJnyTNBN6vSgEdJcSDPpfujn0q314FxM5YyMpSQx9+P047DfJM9Kk9dmPiNa1zO
gXVcAedHQ5DrihiPWZZ78hJBtuPsxKRpN7bxUyOrs/42FZpMEOdR0rQfqko+duMnoJdyHdxAIfVe
XvWuo26b2+bDZPgIdrgR1O3u2hJMMh7wU3R5DSIfRnZdx7QPYyA9QjcAKIIkcz/4Q3M0irx+7azF
bPDlpnfGe8o4e+kCHItG3j8xSy/CWY7F6xTNS/NntETTh7c+0HM6V0p2C/l/qW72bayXasrYwvSp
AalM8hWEXNMpm/QmyUf1kGkvx8M6lB677yiyZ2n5lSHKcO70KOFHJ5RDQIuSwycGu8bztCNoIDgJ
6NkitCBmt7oB13B6Hxjtz4CRQU6/7o36yGvS26yR5o8OEbpnSRBsCcuiwjOywk4NhlzhZJQmVxCk
4kce5zql7/iNWdaz+X4If83soaRJh8NFSw5tYo1vs1PFKjAgRIDl0ly2zvVPvdtSPU1zJ8h85Dg8
nViODtd/s4GlvMyEh+R+J3v6DQ2ZKDalpDB2FsghMvkDwL3muFVFat8ENlHS1yWeG36q38ZrAZb+
b/Ix4LyjZWOxNfjlsoFtwYH9kiMitc6NUTBTf+UaInNmgBB0tER4glLk9TrVJVDb/K6DusYNFRfD
6pJMvwBze7L5MCsYpRaCj5PJ47Jx2FKtrrDzFHf63fLlawbVkAJEOPN1NtnEzWSZLkUOdnw4B4ez
AfsONPkegbupDms1jYb9H4rnQWhsQl5i6Fkqk6PurnEpqQFClsPHLZli2HygBsgDeIeIZLG/P3f5
EUwaJRgU12sybGQJv0jMpSThbnT0Uwr7FqXG9raZESLEWbYX4XeEH+rJZyMmrvbem4eDyA3yELGO
/S0qhHcID0EOS6McVqeeSKTYLOuZxm7lxNtSFiF1pt8juC1hkAfzsbwUxJJVbIcGVO6DaEuOgKCN
ZrvW/nslrZ3512oIHVU2Efs0kwtu1rSeXF/AT4YVB+/YTAa2MVU1mznVxqYSVKFCTP+DZsDBADOl
zrmt6W1JjUh97zQsCyFUWgh8ja7mNfKHABhd1u3sf6F7f/u1z20xr1TDc5tOlC2c+ex0wS58KhDV
tlwO2RIBWkfkvlApqxBbl7Pv3DQufqICXyaaspRZIWRcuYynBjf3LLRTdo5re1S+pcEbmSRyr3Sp
wkkp7G7c3zfAZzyt7P6OA2q7XYcH3sFs6c+s0xuTo4JzhTIH19feu0I3IqZdvIP4TT+P3ExPymaG
AbbeBqM9v9/obwc0u5CUqISQCfeNowfqMy9z2iJRl+sM/5yFN/0s2xJsdFvA35EglyJ2GXbFNvz2
+q0/AkYOiTZ5syGxpAltCa96jSj7Q0Mt2F80JDCQbLVzuemRmbZklvJZUsuIO4m9zWHznNydT4Ys
0f4CBU7plNDoJMwzykkTfA1U40YLSPn9FVy5YUGN+bM3QTOcQRHOqMCjWlEY29ZhzNsNeuIt8g92
aSkRNr8+Y8mv9g12t+KXW5FP1O+EYXYrVXibDNolsi0TW7kGnMHuhDvKLk28CwhEFjYPNeBw2iQ7
lKq1MhcvXZoHO3bqmYqG4EyrYOGjkwpLV7ftw5Iz42Pnpw6BIib/QBuQkVz7MgZbvzeQBr+ui+SE
USioMn78+Jyh5I/Q5ANbyuOye0DWt2LNSHyk2zqhOHkUif8uSJahdVWjoWnN6DMi7LQObdKrTT1v
f+d3hJ04lDI1WmaElZI5a7/g9bAUAV0+P6RVXz4TEG3I7Nt6FoirSfuK+dC96+TdGiEWJpqXLc1a
cSHvE2y5B/Po4ifvjCucVXlCrzvWY2eW4teeBNArUyua2CLnao9LC8USebTZ2ZCukxGesK/ToxBa
f+RkQ2e6wOIP3uLHYMH6vOiwOwyRjQELsJiLI7cPlZWNtSbvFYZrrzAHiZECPyrnZ0am5+R8iJOs
4N6Z2C24xopLS2Rd5+sA1tC3RbchH+RJOwCqybs63oPXl+vbOXTBUOdPTKoeP/6I3+D2cOG9hH+9
X/1g/O7QrI3yRRmZTji2CkpbdbCaJdkA0FDupKeuVz5uVQmgwYX1np3XbwLnalnyD1HeSq+92+Bc
vna2S2u6iOtX2bJCGmFwDE9WXIr1FCn2NvZAK0jKBS9UTM4RA8J+kqdzSEkQxtXfXzM+vAj3RrY7
vbyYaoq+v56pkBgxwI9HocK/B9ygH/uR3UeG2otxYbw9dOhd5sgO1rQ+TiHSBUC3iWbjuyTnxhIj
zhfHXrfFBN72ErDarFoawwz69LeA/kckWN+C56guVRucS/d1ufDg8PsiM6ycEJTpflS+zVV9rBV5
KzohiWFikZyxyHNZBP8G/65eKcrXnhox2gJR7VmGYMqRgh5mw1R/N2ISxgJdDHLjyWsg109rUC8X
ecrUn3VnRMUzI3A2Tp8XqS4W2AG550KlrGj1xTRQu8NOFZe9VGtplmDblJibzAR4Ov2lrqh90lJx
yfUI9u4vQ79mhvkbBELQwyjD+t3sbMg4pbmVNVtmDFsfHbgnTu2xDSCaoEaC0uKoRAMZ5oYicH6D
6NA4r9wMO79SDHUQEIEp/k+lw8eb8fx64qcInClP7QINnoFjanIHvrDc5jMJmNdKux7l7vPpP7UW
y78pNCVlSNWHbKNhqQLZv/ROTt3rCY57r+I+GtwMVfsJtJQZ6/Mjo3A64oYCWhGuVtesm0FoBXD4
gabSa7On18YAoZnbQIbWFiZKLvmJY/66fOkEJGF8bwTC2F63IzqGm17+6op6+6ciZToLDrcHTW77
dZLRlRg7BFFCRvZhgDgWEMCKrrjeljBhTizp7cn+ZYCmC1lW3dDWlyWMC+drcy9RJMbR26j9iFv9
i88fc6ueYNJ2Ju3BXHjQv1IrcM6aM9Jj0wSRB3/dee3z1CQiv4+jyGtfGa9vESMl8c0y82GqOa2N
SehU+X5UqZZZdw2aRVHfb4C3yyoWNhcrOuUDfqcvTl0Tn8CZRyv7qxgOUw6l7OK4UxdBLpXQf2pV
cfoU21I1Pvi0IDH8ZtDjDQGr85+LIF0JhOxDG30e6sV7qIzMyRTC7L5wEpehZg0lmMMHSqU02Fd0
viT0/KFzO1A1XxJgYitfeShzmHcnjCfu5H3edk7mz4taSRzccyLJkLzIcb2xptnwyvQHBaFy4iua
/rTWrHueWT1vfDOAtZUEoFDdEYtlxzvzAOfJMT5xJJeoTf9oWx7XFAG+kXPyu72WU8cDt6SFbQXm
dOUrCfMHpjk0mnGrmmgW0PMOl9Ua3esUh5rdWM2HkUDnTsmSdWdZM2T/w9VXT0kz16M5tZWt43Te
bGka4AzNDe9x2lwwl+Y2nNQU0c+3BikRnKH3r4cnQsGV4zf2it+amxpOQ936ecqu8Z4b+eHWkElj
e6aYC8NcL1fpBzLOTj/WnQO6f/MRXfjHK5bpEl0gGtfSfV1HFBXRKr+3wTDLUykTzafXL8/iXeW2
zgi6+kkzOA28vLU+0WVk25XWeh1GPXiYXU6nR4R3LclBxJkfikpVyuB6udrmYGOYNfoXmURfSg20
4jA2u+es14BPl9FjOzR54wb4z62fb74ygEVKp5R2Jv/W8RiE0eMKUaHfkx7mPTMsPgbOlpMNKsp3
J9Kry571EnuHV5099/uu9wyK63SvM35DLJe6PHt1Fl+n707/w/CP2WKZF/vyUCbdRHxvHSocsHhL
n8QHzzXs4PvhRgcm8i96BpFnN6h3+kqMw8MefZdRy0mRbnl+aNXjMGmxvfnlXHNzCz+CLjyxqKx6
+eAKGejjTEq6LaNH1QVV/UFxH6H1Zh1UXCYSXO5EyD7+ijmI/8Ec+74PXUeYVDJCGy5nb14vxyJy
xdJueAoATnJacp27p5QBC9gpP7cpW5NSrWAreLCocAJ/YUJjYHmDRULia+fQDBtcB80l0fD/QfW9
qicwDpA3UoAZFrm3X6vxGMHjoX00FXLjJLu/8lDMKrtLvuu3KV/HWrdnRDSnIJu9zxsCbGe9pHct
XfntmPNHSkRrSostGFz1BFIGACOE77X1uNvNfN9wYeTXwhs7y9RFi4Nh5RS6IVKOSFY1lRPNN5nW
PbNKSOnfQ9343TgQai7SI+Dxy+UduCFb312oBe5wnL/p0uMiflBeonztvaI1eW9dWo364Hz1u/4F
dUwVNZHD55I6RearQGQVLdlAaFQNrJeqI52Se+fI0dcYLqBT+Rzsgb+B9HZI+dgwwFyl9v3Ok5dq
Jz8YoeM8UiqDSBUdhhwrVaijRGOrie0sqhA/j8OYDZrLryyQ06o+SUjrFh/0+sCp/9/7ysp7VpUU
eEwUzP3UhjfdNor/e2VbIVhYPwgFY3uxEubAuMkF+3lXQVozVAOL5MHnrezGbjdx9IdAHXkTJ0j9
/NYnTZ1QiBCKSgHuI8Sx7MAc7n2OnZ3l4LkKlVEi0373gydb59VvDVXSsvokgzhWrTLVrjDFwJUT
wQya3sbFlxwPgtKSKEEe9Z4Zf8YGwH4JUYjuPiJz0t9s2PAKq/AO5SvOGK4zyvLwB1y1YpiN4Gxf
2ke20JyTZ9v7rc5oUim1Ec8soJAEDUAa0JAJRCfTrbitCu8w8ibtW96h+PbpwUSWwTQRyQGV83Eq
cqyZ3SCnXoxlDjaUOKg6A2A2KaekV1a/Z22/UDlxkBLDkOKYOa8YUjjKDaNqTXSnXRQNcl9SOV77
6cAAJk74gYbPIi6XuxhdWYlYTS/zOmcMZJ11J6pgTKFXe9Q0LLmCxmCmapZhj26CsWV2ZyP7eEQt
3xGSkmonYxYaC7SjOyFxzW5ybjjRjT0uMCH97wSlVnP1bOCizgeNECvuIU2J8OBJlTW25vLycDG4
yJL8HMSOYJGmpsYJXIVzFfFZNnZp7u1jXEh9ZP2bVzscEYMeU+eMa1TZtdKjl884e9+QiGLJ9EJn
anX9RhqMqSR1h2UuPWHn+nwFwR/C2kONDcHmb3lm9b1yshPLgMjc/Bo7+Ha3OW9bzQ8wlO3Z+mjU
rJikqlH5P+REzw5wt83b4rzQn3mKDl7WgwRC5wA5W823lrHOeWJ/YgxQSNWFdrbGmJS3LmodYVUJ
84xurzJWP86n7xuJyRuWogRXQnOdBowI9C9W2enoZ6E6c3Hgnq03+ifI6LJK+p8ba19a+S8EytUv
ft9twizjBNg81uveEEkLLGa8lKklHKgQRWtXkQA907/j1a3MO8eWahYGNcioTkc6s8lyREO7tlxL
u+Wi3UsJB5+KBO2siq4ycUo2RduabpPIF6BmQsUKLGZSdTbyiAsMStTDjeCPz0JZyPjDreGmSy5v
n5W5h3rVJ+6jVdkemAbHvWfGe1vqu6+2nA63/2dC4GW2sCQQrReqytxgrylLXw2rQR9hSosPRP7X
J+4/BQ0QXnHSDV520nCIE9xgW29eUS1REsc8afoZt6AglSKbi41lI/eaCEjb3r9XlU0M04Diec9m
naYFBIRhHcL74gFsnRvwEsAhd2k259NPK9BZcS4vnZRJ+fgjw5szuhE2r0BXzMbn9BDDwW3+H2I1
bN75c49MPRBHdMkAugt8YZjJQYlc6espSRKi2xCXkR7ffs15KpubQ8nr/dT4M0QV0nJdky2lC4Rx
icXXy9aGpcCbHOIomMKxppEr2Ke5QXuVshyuuNzM9UxfjNuqjjTrlxGq2zJZqVIF9mfQIm/IjuOB
Ld8dG9G/BHAdHniil40VRO/iwwrh2HIyvrSogI92NIWiGNKYrDzgF72U3RqUzKk5jrhh6grqQlxF
AG4A0KNMoDP11zz3NbTYYmu2V09zA7MMcP/j4Snb/DYl02UWoA6kZm4E4tpkh3yLe9dUHt6MmdQL
cbo6ROar/+O5lLC75q1uatsbsJnonlsR1dOcTtHLVv30psn5SZjpuwAUp6YoOKbBXlj8LpiLR+Bf
O5vwJwfvbB3/TMUmh2kSAM7rGeiViH6sWHNeiuu78m99kJNUb2yk6vf940iwwot/gCtZIBNhLpo1
cZsOf4f4vNR/BXAhujmKalYmR8thp3PumbJD7f2XbWOgbEFS7fnCSvwh+svPvi63XLAiLjn2yAnR
HDPND5c+dCTa2gbQzHNOE0pJDXmx9oBftqqWcybFh1844bIpw8Co9sZlW1IuvtfWpAaW1IoRZjnM
TQlK7TURdsfgfxrYbvVzbCrcqptqmFniewNRUNyXd5zXAJrpdACGEXD1PISUq/1btR6JG7kymQF5
1G4F1JPZypLIZd3FCqEl63HINuPodkOP5KhPkYN61D4po35n+koCR0JTvOyOCwNfs/q6jzy7q9MS
EHDph8CXRtUFd6ZbuEK9B6gyQgQz3+5qIOIIOgSGm+HcDr/ltG2XtlRGgq1AVTH5TTmEgXBb1kAC
l1h/fShMC+4X1aGkMY6p/6cDy3jXb3tNWnU7PH2PUa6122FFQ6uADfAmjVfmb69+5sWrugBba2En
sFkbGDl6sez9rFV7p/SgZGSjgarYOMRWzKlwVQ8PTIkzBsG94xBbYqVP+S/lDFWsBeYNqdwYWfxp
cu14YijFMsu8TyQlPUbRfnrzUo9KX+vRR29wJ82NvYpLrlAMitMpODYnEWANggQEtQFyMUO8ka6H
z9+PJL8Y6Qapsfa0M5ScVEzDSCf6BQWljUQWVohcCbDMOalNnRI4sbiSMPMWw0ubH+VvHaBYJ/3c
Z2OsdhB5RAZyKMxAOyPyM1l3AxJLlfhxti0SqVZ4+6BLW31sKaDo5tyFhsemXWcQGbDsf0tbhzGt
BuOrogpaW+6uIcaeDWPP/hCAVfileqBNQFi6Kde51/u4X1yvk1TKaMm2xHho9xNUiMzSUDVGiLDo
gLi3piqJVqkXzyBVgOJV1SCY5GvYU6VxEpSzBjVyP0czygeQbGczAy1MeDMKwvdktIVdT4AoW5Lo
QgxqKsXez+531rsu6PU3wMk6LqwgDSoX+F3knX0blCgE/2kU8RSJXNq0l9fRX7bfNz//hdDIrkfT
PKheD56ja75a6FHvqJuN3tPAd82bULU9IrMPfkY6FbxVXecd1VazWdIr1Gj5ZCbRelzGerczA7Yh
JtPVbpifZDbFu+I2AVHb08x1X4Uk2Le/r5Cx95XJ44cPJDhgfcH4iqWorrLJLPFDozkLwGWTn4nO
Vjp6rJ5CGLLliSErRQyBTXY9H7JNA9gf+B9NEc1xHEwBW+xODySlz5E2rsz2lGhUYUiSg8DAIG3U
AHG1bfSvtM6QW0Ewbn4Zc2MvQDW+QVHBmTtsuLw/dW2dawumbob3NSZaDlJ78ANdbo+AvNnX0RwR
wSA40PLC1lVuSOtkFENOb/QfOtU8P+AoEu/HJp7mlN/bLIXraKCX28F9WkwZmLZPqQ/DMOvzC+O5
58UgrJ8JkqZn7XHd7kUGSmGdhOLHMidyKykPL6EBnEkrGOQJbrGStszwVKBmA7UTi2xNa3R3vrdD
+HA+jbk0IFc+ZLAq0PFVS+6objc24WdUXxKDu1tBJ7DYGojIzbZlHiuu3VWivz9Fg+F5v/Hk52vP
iS8VH2qK89/5JQwDaJTQevkpa+3ZBwgvSHo+CDj3w86eUS9tH77zmOKmTh6iG20A7tQw6YbEyMZ9
vVgloNG4MWxNpPM9UUzorkYQ6+j/fktDzBZNFPXnRDVs+ajKSJHL36HDAu6KTRnW1X31WyPTLsGd
MdMdBFnk5WOSUdpxs4kcbfp4AkzSO1lymRkrvK6Q3Tj52UqPKNLfyl7JhpM6vmoK41Gsg74YkHdU
np+FSLo3FphocA8uBNzNp7B3k+MpJ5QV9sRBP6vyAOo6DD+KJtqU0iilTWm//618hSb/XJ3/Wxbe
YKF+TdHMpH537KRxEnCnyNYivVdeX35u6C4zGcvx32mSgNJ6khluIuSzCeNvMMS93DCbrUmGxJFk
xd2BPNl9eyW5TwlY8suRXBc4mSs5vmLQtJKkQAaOKokDtDYggoTDWHbXDtvHO+izpE7V/Lz2y6Ez
l9N0zSHsnjI74A1mX7h7HRWz6y05UVpc4Kt3yY/Uv0BkDiRy+U4FKqNAOLkHcbVVar93nXRTf8ZZ
dl/z53owOx56HYF5gL8LFlYn8UpBUAaPGV+5wAWD0p/0laEfVQy4viNvuIXsoXEG5FXBhkOtQDj2
Vdtcw6Xk/fNbl13pW9cpUe1qIKgVPW4DR3bdhXBUnrCAZJ0Vz60JuOigfel7EfPNMbM9m6GAEYV0
nOI9lJTDnfR9fiEzwP2IxCGI2fRSxYvB25PerZLEjIdXYCuAvqqxOF5Qsn6NbladAGpAddfZet+u
obj1NDJCFyl3oO1tlfu7T40m3m0TB4YDU/UtqDAnI5SHCXX+6VciZ/Dw6ze6qgAgED5fi/rbIj0l
qPfLCijPNz2m8Lq/Tr8fPlVvcWcGYXtCaN8lEOVFCvBzIqlN8c9gMONWiVwxekmW9ifmcHkNPjJ/
IvDDgJ3+5PYlVNy8yvuSs9MXZ7p//WOqkWLUAB3W/2A+JR2jqE3N4WSEqf4z+1Cv15g4g6Wox0Cs
xaxA5rL/i7r6+nKwKHWMUmEazsFqJCVbmUb8UsIoVyBUBr4P6Oj+ob7LN/FOSqr0uU7ZUQ9H8Vrz
wYdic6l/PZfwGpjJp9Aen6ou5bFKH990UB3OusD08PT5wnzxwhu7/cjbxHTUdXfBQWP6x6XCCqI/
6ATkBKiA6x43Lo+3og8qy3/b5xvFIIZbzAqiKYvQ5k7HCd+Xbapfdoz69e3fHlkbrbtGO5hW3GNl
xx1XZ8GlcmGDz66z9tle9aNr1Yi/DFclBiTS5dFRHIHhCMnJLEUobP4okY8wCj5/oIyy8wUGm+ea
AVWTAzhkU36oP4CXWqP6zcxmuE5SpDMg/xxVxZg8/fQOqX/lDcnd+YhmC21LaZf4IoNeoct9IX6/
i8H/tvmPLcQSZQilSx7iFo6YaY+FnpegOI3kwL1VokUvwMPT58XyT5BWX+WsmISvy7BMY+MvxR66
jQb4HsAcgourAdLAQ6/FzAQaEPFITgW7llm7D2+OYq4of1aG2LAizny5JjtrRBwVrpLEmmaJQ6cR
sUhs5Qu8sd0V3QWjHlILs5CAg59SLlqKWRcqragU2B9/CerxEBNf+a64IWFf39UzRdDxG0WHz1So
xjjor+9ZcP++MdPwmNXIGgrrbTzkd6Dp6M3ikwdG4oXFANWME7pHzPTciCSnmIxqV+qy9SF1Ods1
RJxezJrDT+5k/B8ueA1mQpeF0ncRQkHvpL/P4teWADxfUkLHmtLObz9h/um/X40S9mD0eHOaM4/o
HI5+bagDfetjELGKlI4f/yUUSf+sckCG4zrllbEYFcB4KQxczXx+Opl0boTE5eMEASkUEDJFKe7l
U0ZW07aBvOAf+JWHCGW8IQ36un0hRmWqXQqxp0hgc2Pt8xXTay2YVGnbplgNylEXPZlLJvor2KDH
BW4mxGUcvB82rHxXlZ3r2OfjQIhrNSxlt7CTXV59q1DXTBwsuSBe7m3RHN2OKZ/nZ8VQwhAB/2dT
A1Xg8UulOekpvwmOj/eAwytg6tgyRur+nCDQcudAwhksdgKUiuVG9U1R0S90KOhOxmHHCjC79mR4
cH/xsGYcV2DNbn6RRCmqfrv/mQvzan1pbBZKxfS7dhX5WIXabq5WQoFY4pVxu9ZT709QFKrE08rk
4pyhXpc0WHaAZO8i5UKpS2+Z+BiRMj2h8WgpCpuOdRPigN8FJ8c7NdQxJWj7iiDKraBO8sUkZuR2
wInkEvcTb3OP12LkleVZ7DI+jEgIcin6fVxl9gChsHAciimWW7D7oZa23a+/V9yf2TSfZjn1nBPs
vmgIjjhxUl5tqxHnxc7Jd9Q9zU8qnxICRM8OVGWoSAS7W8m/iUAarstVPNryOf1CZM7REro58MWO
dwSaxZMEfCExw14Sk2ojOI4Pl9/D3FwZv6porraFymFEJDUMzG5rFnzMVDLhfLtjTl+Rz2DeDvVU
OuBs/mrxINsoA7izmjOao7vsJOHRS4GSR6oNAITXQMqWxCNtDOsooxh/9q+KIh6o3RWY+2kigQsB
dQmqRcqHjlZpEhwIkYfSgxBiijCOutr1IZ1+/nbenTGnJpMZuR52NQTOHi6QvZDivhnagH8CzUQY
qFDKeYcMsi3Vo/hFDbefZLiKYcDpEBm2nXe3LldRGJJmr72SZHAHq51IgMUoYOBA3Z4J77cwSTQ/
wicOkYdbHcj2jxAKVN/euYOywOJ8Hcrv1wlfdC2iDnbJynZeaKK2ywsywy5SAzYinhQL7MDO5zgR
xxqFSnrpqyRG3z5uHHqHJ9EMtpk7in360gOLxogH7uihdtvLVdt6+6mk54G3ArnrQqe09i3jsr3M
Cjl9KoBPypuP/OcRa3RAx1R2OD0oI/vckaAZkjGsLknbRsTpN824F5a22T8XPFN13jUjenEyj2E+
p/7KiQX9p07UPXMdhMNvEamTSb8YQ7DScIfnrHSIqe216flfx+v+JlLqcw3ndxlj5SKB7hm4WF0e
Dc7ihQzWWFk1TKK6ZssnKMJk5ufZrWSJ0zdhLjMZJYOHOH7H7Y9P8EbDt9q6U0fU39wWEQC+JNDc
rEwc4m4gAYok5k5hkaKiyApOujlfL904OCsGqN3coyE8yR/VTssA4ZoAIMJI7mFf/tlAmuW2xDdX
0Av+2CVvK+ExmNzg9Gnos/BTwXVddwMgVPjBPQ0SPvsjPtkGY4mLgfFdNtMF15YQ14L/O4F2BSk/
EyNrW0s/CxXgXLcAosy3Ewe3K+Otn0xBy3/CeaJReFcjGOTOoFbuuxeqyVYPnpyT42Jd4lPgVeLm
ETZPVhi3Aa3Wo9KjtsPIy5fMphSDGtPH3NYPenF0bfNa8k5BFUNxjducOlr0ue6yNmcVM42G9kv1
2DjvM7soSwnQr/vd8T+PDE70xQRLb14VkqBOfYU565r4FpjWy/OhkRZHG+Lwmpuko9ZYzyh0RIgd
6bSCoLCjVtZAPSusqjH1RVTEADr2hZy7PMvMFnUM6PgCi/BWy1wjD02vR8PLWyRVLZK0+79GbCIO
EQscWKHqBohQWNeH7T9slQ4foA7EG0gxIOBbqRxl0o9efBgPoX6v2LEEbTI57wYBhEbPxSP0r0Jt
JkZB7kUtqPJPu8mmN7HXbeHk59zapcSm72L9ushIF5NO8S930HdKUdTDsPefuQkaYMPE15MtJyX8
dcJMTE+UfytEcr10rQSgla/mPh3P05oFZIJQNYBTnFicoWqzO8UG9YQgGkq6e/aJ/+Rdnpp73tmd
GxKQ8d+/oaBxvL3FeEU2QfhZzMVLJ78uZuSQ7OSIQGTpc/MxP9Pf0avUZFwpSfHYWft+k4szNIWN
Sh99cplDqY2pYiORFRHaeRYmJ83u4bUse67kmA5Q2PaByEUkUvu6mv/23HEi1wJlLdGyRjeZKWhJ
B2rw3YslyI0ilmvC71jg+QSbixThzZJLnjN0xWsAFFTGHEhOPvJRdOg22ptm7cVKPuIyNFzzFmat
/cADO9UeYrYl27rCXfXXVz88lp6WYHAglbo+sXp93iRjENEwhYLxw5ebwsRhQGhEpk+Jb5auqxOl
Jq3T1KajAWDKewTSyG94/AFUDHFRN6k2lH5I0UzLH2w1Dl81KbmGQCaDKTFhMxlmlGfh721VdJXW
CJliok4/yBYURBFB5pcexxkRU5P5c9b1eT6pc8RZ1LrJHaVPKQE9bhUzqPd6VY8jR3U97HijEjIv
2bpz29tTLx5MaR9k2I9dcPwLNeJHh2F4FEO4WeJc7TusBV2ZoWJ43KxP3PkrE3mOVtIV+I3+2HoK
Qj//+TsUbu6RjFrfaBHKF9qxT33edlS1f7IH19FO1SL17tXYACOxTia5FkLQQuhvFnXPD7J9bOXB
qvspiNtzqMPkezPyvScM+s43abJIsraoqnqYXnk+cKUY4qGvWO5YaHL9MX4ERCVJ18XmAX/YUWF4
7S0gbB0WOTjohplYD0DtwxHpRl405i+USv/dKAyc4nbIKsyp+PSaDG6KCJezmG3cOA8Ucw4kGizT
sCUQN/h8XSZROzPs2Sbo6uiYCJt2RdH9A588C4DO5DTXvcaYYRjDqUqC2J0+YgywOkSso6RHHgqs
0+uf83HS7oq7JvelWFwoQdwV1SfZ2l3zX/5HprkD0Yq+JIW8zlsnS5Nmwz4RX6NShRlt2IrcKEam
t1sskF8OOMjUs5LhbKRnXiUI9NPMl1pndwYEApjiL9rxTiQ43UJeus44DFc8sQBMMl8nK3d+6kRI
rQxkzwbcYFod3M8n57DDA3sXHSu3reL7rmo/bMLgD8eNlr2DsZvBaXbEU+r1Z6C4Mb/Da/Ep4/9J
L3f3VeSC8cBwT9vMJP3kPCgSC9NNMWuY0D2cMWkTBcbt4stv+an/NYFjW/8eEC8Sxk6vUdEAUclr
OPOS0ppT3Jidbrfd7bTYeAg2JcuuPO4gK+ZBNttRwpkIlhstai2v/9xlBzPPsK6yCFOzQGgkc3cd
LP8zlLwJ3TMcb0ap0s0s/lEuvUxGOzeie6qwQIX7vVCGUq+sk9HkrDhG9oPufBNSQgJ6SyopTQAC
Z5wK+8UGp2SQR7GuZWJclTQ+UuWcu6DSQdWYCUujwQQXzCVDOsXRcnFHAZVfUBrPc13eqwy3pIkt
J7quZFoYrFBeXZIu3EYjPa0lKrLTYVmVTJ/Bj2dobkEpPTibAcExV2MRQMvoMFAC24GIhx5rfS5F
ptMobAdJnwR63g23qON/w9ZoubVBLgQyOjEhTKbzjOYe9N8/6qFCGD2y7vBFvzBSgDkCmnUgtv5+
lM0SS3ew9V4nChm39DRy376SGX/8ihZL/QSRmrVlZXvVGf9VZQPsupdJUb4Ye4p8G2p3sMfEox/e
q8LF1/ShJu/HOoG0G6IYAwwnHBEqXhlNOB3V5gcxB074+kA3DPcHgJYRocaKjQqEj4vDNGsr5WzA
5qJO602uEDPL4JLPbS+X7PgG13X7UqBJxETnhdrBKvz7kHoVn3M9WEVbs5XzHHaCn43k5LWSkLlI
n3/N8sg4eU3mIjVB2sFLH+1p78SFWFZSYFOf93Ahs7O7HJEf9SxUlWUK24PFuSVhdtXE700agr3T
dysbYWaLw6i0lNX5Wt3RNq6lI56A9yhHUhIDpm5RsD94AtAl9YTjd1iQHcJDOUIgwhP5ICe65nf6
sBRfYY8YZY5IdL2Op5OuUdxZD1qBmid5re7S4Sv7YGJcd7VJO31oXxDHNWG2H75pZx0gGKXX1UPV
wmQ647YKqKJ5v3zX5HKEwbGW7iQY3nHGGDEmaXCOL8Tt/zWX5FwV5kyPuIn1ClvquLDsr1NjgJvL
o/UypY21xsW8Nqv9vej4mj3tIIF1eVIjGUw//l13THnZ8ZmO8cPPLh1X6P2HdyuJN3OBZ9IpP4gZ
HJOOuFppvMZMTPtN8MKWIFrVjFvMw4Lb9dWtVw4rFT4QA+XIqEVELN4FLAbdvtJ/G0AP+pFhqDpx
UtHTnGp5AVMHcN6zjLAZFWr+iS1fV3Ei3ZGcctPm5kHJtwyyhHZB8qXyG8v7LCkXs8dn3Kp42huY
gJ1fyzMY0H8NYBwVFsQc9OJNiV+bqD+mijEMNXqPMRLq/Lh9t7nBz01fS/xCBnjT+LnHuq8LMnue
9mkxcIzvkm+sbGh6nFyTvWlniWQJHNYLRSLIYNbOzrEz9+fZ254DIlnA8PVeYM5gMnv1dkqRIGOX
R5GO8yayRdA48Xe7zKVVy9Sl9l4KlydpFLPOud5KRmEnDfowh5je/RwbzoUrk18RlmxOPUFXOWbf
ObW1qEPjA/risnhQeG9TgU1j94X/xS6z7JLFCjWdndEQNhKjHAzZahOeOsdDw9tIzAIt2qSB0/Mx
YHIdX65T9tNekeTzi8WwXO9nzswPcx2b44iDwHMHGUY2StvVvl4+muooHlk3JcpGm6Et53da/Wt9
Q/K7hsNkpv0MhIi528TjrIE+vix0dwuVKzhFqh/LsVLj9n5VR3xjM9x/HiwbrRK6extVeMSfy6XQ
t5f+zwOlI/BjWoJdZG49/6+1VCOITHK5DeREodC0JM29OlJ+t/kdg6fLS2X/HHBx1gbnC7geKdCh
hpxvI9VK3RDgMSUajqlp/nG/hGdLkKmy+fyUt3CGWGpvaihuOh6kt0o5SGYpzPZnsJNm9fQGqQ6L
pDB/BIRLQsO4RzNzJoo2B9h8fXU9dYYzdqjp0/z202mEAiXD1bVEdgIypu8UNvMY/j2me+aSiS0f
WGLxWexqzgdKl1Vy9LPHet6EkslIMalK6NEeB6H62g7BGSw8ADaZqlyzoEUbzy4f5ydnQHZtD9Xf
udhWIN/JNIQ8xW13TkdzbcEp0I23wThH8e53wR0UjUWX0CfmpWvxQPVZ6tO8UsZli0SzMD8zqzSF
qJjI+9E14WGxM9IF7O+E9HNTwfd3ikluh2fzgYs55NkT8uSyNfE1jmia2JKYp42knu5pKJbNP0xY
Myn0DelOCYur/nEBK1W7JB4JLFXThO8wRvLx3Gvd8ELd4cYbZ8gcFMg+F7k3E8jkclsovrzpIihz
12MTJzuwRJV38R4zZlmfxepp5szlRcs7YDYdw8Cr0Xws7b/uiXiqHckDt+M3ynW0cfW6LrdhlWbK
VVoTplw0qzz3mGNoYvzVgKCiAdCy6s2P1fAoWxww+MKxY1UiVwNbX+16kJBUtw51KfQlefurjThB
gxLusfV5sPt2UcCtkElMGOqZVdAZydexur8xsXggVuBcSSf/vOrDunaf0C0F6ULTScqGNyR6JJ20
Uyt/oUIOCeH80nXTnvQB2M6ayozG0zCrDCQ0pZ0XBcwI8XU4tr3fDdAeAnCE2ulTaBa+BU3Y3Fcu
kcx4j0tdJozWoOQehuzePcj0xmWi8H8fV+bQWqVWKejKAI01a/MqqSe162yax4SMkcds6qO3S6i3
/g5uZWaigWqvS2w9LxYxfYd3DIequG0F5A2NjJa06evqYWdt273kUH+pyOLVh9oK8pE3kAO9yBxj
GgXWXPVHfGd5L5bFWwmMS58R3nv6DLazW2bIs8laQtj6sV5OkD6WkR0tqLpvgvYjnA6bRULNnDNP
O8zscN4nhS7AD0yQyyKyNOjJegGw7eLt9RSUggvAgljC4BhqAAyf/9rFShTcvaT1JO1wr1gssEVe
2Uy0hqvM3XZ6B6IqrQHuyO8RI9re5Asl0ulIfwC13uq5a0nHbHN63IC3yXe/tQQYacBGgO9BHx6p
LB9Ikr+6GUBLHaw7tB+2fljhxjQStp+b224IvIPSfvse2m4vgaOl6UJTcNvf06ohwKOD/7I5Cs67
t83cwYebONZYhO6DoIju6qx+oZYwQXKIeH48PWrXVkG+qMTNeXHC4m5QY60x9jMsRJmPJylzobrK
yjSpYkSbs1Vz0wADryzvlcBqgJ+w/STHdSUN2IVJA5iwTpA+QpOl133oWU8LC9aI5iV+bqF6bsVA
8lqVy36xxdOcHE62PBWH05xQNUFz+kJkSDwqFWwReCpfOJx8ujEQvgo91NLvjSdm29fjp57qE2Vk
DFb7FuL2lB/FxUC27Ea/9NKG4bPMvu3mkeRjPFzU5J+Insz6oXqEJhR2FncTFZT3bztpzcf+YA2J
bmLfInuTTKcF/EujsSnbSyIaaRKFshtCEIgbYOrhl8Q6LrbCFGK/XlwdFQ0RSaEOYNfIE+vSmjfG
KuXQnFOTKWq+SNNeCTFU4iI+q6fJrKHYX9duUhZ0Oi65OcVwuIj1fFVRD7oRe7rmhUGysndX5AYu
3vfCjywC+WGwj6pAdParJbVI5ikXVsJ3qMHO6D96GnCIKw4bLmzLzlUbvwe1xSAWwJ4A7w6yqJCo
rqhS2Mf37kVvDgYQx6TRimjpfDktF0I+YYpztTQstFBifvp4tdRcPNXWpGZLg5IIrI0O9qg05x4e
/dYwiEUaS//XU+uplq/WN+G12I0KOiqyZyfYtA9FDWLXrl8yxCTzven+ZnmYZwKi/PSLybENSuUN
K8VTBOisFUbfqAtl4wlz3T8SEvUf5GT1zkKinOKlVQDtd7lUU1AkBl/8/LGS56Rn/7IM4kUPr2e3
KzU2I/roQe43wpteSweRMQYEP/pr1PGgvHox2gnVtRrFRUTzTdR+o1v5DVb/2t+RnYTdc3PqrTVV
ZZ02MW9IMzDXVawvrZ4OTnCPny/fB5y4JIytsbQFD5y7JGVwle7KSeay2VDzkPIueJrIk8poe1Ly
ex6Aux3Veg7WwwOzfYT23aay3d0WI/2rXQC6vWHNYRZ4v+LXtwlDamdZB7B75Kc3fPQ+iyqT10zq
NF7oGOU5Um/XyytYwHVaXhJHKZjln6JflRaaMETDPEA/1b+lO1xDiHXhDoJNRA3ZqTOi/3n0GA4P
Wof8IPy4PLn5YeJUtXw698PmH+OcrZOSHFfD13AWeVHKoXmps27XXv+7djU47NLUxmGTTzUc1Stv
7piz93qyfueihdhTM3J1idZYUQbxpwaf7mH/eAqbid84f1EL2qsJL/cMU+T8wrZeAgflM21srWkr
FG94sNJ0xRmWwA0WpwGLjNuLzkNeSLn94V/GXzgc3kGG6v//3Dx6CPb+UcUkSrW4bZQ9ikU9gIVT
zQ2oiNZgRdNglBaDG918BIa94EGBWwtYT91LTtg6v3XRzZzfRVX7HO8TGMBjRlpK/4VAQ0B1HmN1
ndJCLXZMDpA3ziSrN31x+GDxwwmcDA3CqFgaZOAgByNCnji8JcQbJGa0BajNtqWfueGbWQt50WSz
pnmaC6SFIvm2lM1wE4C8KOQ0w0IEd6mgOsbRSXX01j84q3xfxq4kxDIPzBa/AFj1MA33tPta3gPb
G5x8qILMnpxGe5vErzAKnt6ibgmqoIOYzkUgjUC6WmyHnlA358l4BJAWUVPEHmb+i96aq6O3QVj/
bOXUE6zQb/qREg3wQZD53tKHptXGLPYXF1gQ+JeJCcCNtaRkTUpF5mBvZosltjNgZ94Gud4lfoN3
H1r/pzQ/NEK9Jq3DQuR2dvl0S9WMU0ACXkbdLl2HJQkjJR48RxtYtlgh6IgqThPvOs2W8pdEUlBo
YLfoSePA++gHFEc8wB6ce+ik1DRgmUN5RYs6vA475ujLP56gxc4Fw4TzvwV8kA2do/7j4kiU5DxN
AMO7hfo1FF1IlkB66qaXYv0aRc6tLOfhgMLSHJQnUe+t5DWQ0cNo4KLWhnUXTaUk2tOezqpuodYj
zqNGK6IFsNAOmAM0QE2MNwaicxxwRcoRIatigAT0XmuOi/cn0Ej77Rp6R3HGFEyx0ekTaXx9rebd
2iTW/1fH5YS3o/n0QKgIqJdylZvFtfjfGvXfp+xNd7zgXY3vz0U2vYf2AUmTSciuVL5z9tv9y4zf
JbYNYTibee8mppIQp2Cp8LrGbvAB35R8pXF/piBopwo5rOd7rP5UGbzia7xcVKlc7lLlTaVopInz
6yT4YyuwAoPXP1nbz88+L5yAdA0k+KoJiYH7CWh/hP+Y9f8Q6KqyeZkfsM9uSWtNdQcHBlqSgerZ
jMbmJtBRjIn2MO3VqKCy3KH8ubYRiMzSCr8aYLSPpv4vUsL4FozF6mHv9++l4hLDXf8kgkLM0Jo3
6TEBts02eyD+tBEcOuVtDftBnSHcjXkiDRNu+USsG52AwBm42+ygN/rrxB3rd6DRHdNuewg36+EZ
spoLcW7We6BVSxs3Ss332xeF6icVQu9QehUrnF2DklL9stwJPabPQoHDyPxfaeSDdMzI2fYx8SRP
6k5Xab7gbD3trQ7lL+2wSu3Smay94iO527B/rj7q5waLHph394H/0G80mW1QLfG8+D5watCvMcov
fNAB8+kLW5C8nCo+9GVRnl9Qwvwhw/csr423FqfVoom3PS0ycmb+0oNBqTqzrxt75aMzS3rEdKRm
THKQOxZ0ro2EbeDa2cmsZPf7yQFCOUO9Yf5iW/iFVHEJaNWFa0hsUY5Vj07yNfR6TuyUQCJeF8fK
eX6TuTFL5rOzpje5Xh/H68UjTbE26QfJySeR8nkZh62xieaZerFwFHth2MmgI+tpAC8GirNJ/yvF
Bu84Gxfn/X/PKOUcc6FPgwYbXdBv7N7UIeufFBaTaVwp+NLFsfqhLliF1Sn1f/fXtlHsVbH9F4Sp
uaUwRzPCUccvifAQPeVBjdiLf6pxD+Nj6jYhWQShafYAxMcC36k5XVD1j/2NB9XAl3eYF+CB2n9r
hw4lnsGKGx8istoONoHCMAtWAIlKsYG8y2mMBT4DFQNDPMRmX+8fu2Ow41dlbio2/62qYxH+qu4N
r2w5FexPuezh9KFaVyzzywckKMPtaAeNA8gVODFKFUN/yPyEWvcW1eJ2qBHjk+gs1WVwWpaRprm8
jetRNClonmWhd+HP6Gp70mIj3rtrz2yH8QHfZ4gy4lxHs0s3eNGUTFGk2QyApUsIuEVkma7uVa3I
YhK/u4Oi1jsEpL9W1cSDaui9tn09yJ6UaGXwLGhW6u3WrX+RPWjdn40N1cT38G4s2curzGbNPF2K
ZExsOBrkpMwEvUdvNgMEo2yE0NJTM0jskPC7nZ/8K7MvAVaGhuorErLoaZUpHp0oUMazcKjl+1RB
54ERa4AIQgrDzrQzOq4yK5BOJW6FT6X43U+cQYxMqrwcUADdWHtlgtLvN27YiZw+cm3IVUHapaoC
5v36zceotl6AGPcgRKiDCrbmViBlG1EY+po5B/t6+b2jKYn0uIIt8Ga3bSZ+rQeosQX+Dmx9GRd0
4HOtB5wikxYFcofDROY+zurkD2K3tqV+lYdUcyKuLpDhs8mZm/RyvAh8wM59aPAr8UnNbZnM06TD
ZF2j+e2nhTH0FnoQUcHP7zfyL5fHbA2Cd1VceylZHp9c4br6RwIm6s5drODiNdghNs6KPn/wRDi4
3p+gnufKI2KVy2izzBAKslAova9y3P2P/+C6TGde6Fm1t+YYlIk0Kp9tVp2MfweDdZmAHedejm87
HiwW/hjoQLMxZ6kKwMzsmO0MyohHUPVNgklWMNyvOrK6rhwCwwFeaAWkm0x1E66pK0eUE1s3iFj9
zXx+ssDLR6AEDSXygMsmAO1+YHCrAUf2qfLUGnFMudU7KOEHrSjyC3nNo/gPWWPQ5/QnZBUF2Yo1
PMxBJ9rAx3tcg+XNoQnzTIiKrre8MHqYPsS+ekcmC9sVtRC6/QSYLXh2D8Dmo2nn8WMZdmqigsO+
PId5UketUQOCKknd6bdHcXJVWItM56M0vdjD0Qz/afTgOtZJbkjlENv1aZowep36MWXqB+Vg5nRb
3HGZzUUHheLZdXzLn+WKW/vWVq8jz9pc/I6fwEt23TGGqxgnUGYF/xFQJ1JW/SArz2xXdzvZneZl
D8UCggCb4ZrVr1s1CU48ruBDlCrGNe7CtzIcZJIy0OYU6mY0Xls6c8YOgmt+RfHwA8wEsUGE/GC1
n+h+fp2uOJNllw5jedYmFVZ3lc/ozDO6ZmGMRxySKMUvZTsbkvXTm4YE43JXOCYXjVt8tSAt9JXa
qkXfEefjX9wOO4aSAffoSJh0uUnwVxhH9Jb5zhdvlgGET4y5jhjAWO3c1++iNC8PGMO0nlI9kIBY
V8fIl+ex/yIRyp+4YsgV2XwB+tdE+pOtyqACP27JrZwt06TpIuArbozGlUfYXuoGI3IZUJxHSTAw
THFHwbdw7ixQAyBWiDWhhvopls2e2oBwLqRy/3vn6GDleqikKI7uERdlySe8iWWrRllVhUjHLQI2
ty9uFFGxmXdHNwjS8u9pjNQyaQBIp8RBlze4BLI6iH4gh/xPmNl2fI/7vZKzG/24dPk2aprthsuy
cIrAVcxVngh4jmQbVGhp8y85BzKOoo0T17W/hLxu3gJYAHVZKL9D/bY4OzWU1TrkDwxvPUg3umSJ
KPQ0LPzolvk73yC+fq8wfb+4kdupHVEljjuZUmPaliwaGeYdmPHcYo5ABnuMWSWEYJd9HAxRux6h
9lHssZ+lIpctbDYwTKbOWxi6tun7doZ/NTfR+kj/ktTnqUh866hAap+wx/9tOOoR75ss+kR6uJIY
xQ4aXMfD6wAP1m8iQrM86cPJVF8SyaTxgzM+Zaa0quD9wk92R5jUaLQQxclCb/jrE1+tVr9Sbk/m
fOjPbN2Xpj9UvGpdXUGkJwAFxTMlwQ2jN8qk2iEZKyAZR/lytK5jg59uKZuH081jjtrUvCk2B9oM
JKptO6R9FGTSag6RN9RpBN5UPyqSUimnyV+gSGbMhT07TfhhYT2YeN+ZkdYw1mLZq9E65+lv+lBn
VLTbHfjIuDzofaAHtRUdxq7WFnVFOtHDuFVWgrItLl6QwfbIlGgIsY7PKWH7WwPHrEWrJwz4sH53
uxNIqOtNWg2AVHB/gqscHaXmSF3q5Ove3hPA/TzajRwQ02cwxNhc8dll2teHxsWFBDXUkuB1Az+B
cxhOEK+p+XVqJ/3ttVv2oP2wkVx4anmrlJkgyGtnLXxzLFceb54RDUKESHBRDN6SAFzZAdbAMJ53
RfCot88blWgQZJoW31J+coKd4+Q8cKe0CpJ4J3iCsKUJLLKTtbiVbHUn+D6dugrZDjSqjkTE25/F
lm9kaZszfeeWB63uIwHsJO5l3DxKeY1qLZsh9bS8Uzxu5E4nsqzxQbL/1l8d6Y3jeWoOrpnoKXs7
1tzpWEG7Rh5VX1h9lJh2Ti0e33oFqlWUVkFqxTMoSIe4GbbYZegVQaGU+Qd1jOoV04ZyYsEGOZ53
Cvee+PLzADWXqf+qOpy+HENUxdz2/FkJ560kmOjijp55DqWRANNUaSfJcGc6JOgksWT/qZnIVmAH
h1ivJOyaM4qP4uN1Ib3ZARvZhaGkN2+M9ZsM8S5uHQ/zquEUM6O3SQRH6gm/fGEobgWlJCLxhZn7
oWoMhQKLaj9UNHOvHswVhQiOXozTlwbCB3mbpJ/1idLiuzMbf7/OEC0hORt0MbiSLW/B9T+Uqj9L
JX4qHK7KmbvBRIYAzWyOlSsBQ4RuGo8dG9KlxRRDn9f3yngFCkMXjw8PI5+gdJ9xEPtFh9SHZK0H
i2e7ideq7rx/6/pLKx+ZZ2WNMBYbrk70WzekKFk90Y1OhqK8P79XA69p52ZRB7n8LmNLGkaxblnz
9/lL6n4jQD+scI6a20Gb/l8wUNLsYmFrlDHCUtWiHAhnImqRnxOsTgtbaypq16AOFLzQEVaELIAQ
1YXd+ZDPfcTs/MhsUjeVx8VedRMuE6+whP7z7Pe5m+WN/8LY+WPns7WrBJaIp2tLSX148oUFKvPB
aUp+RiZj1afd+03MfWdBV27OQAirXhWjjpNfZN+ZYAbnneUb7lPsqE1mPR+qNl3btnxD2pboH5BS
Bqgitb26oj9GihvQ/oFNei+szjr7fjDbLixEm0OAmbGyVHe1YTd34peium+F13SvxW4FWCpG0Kuv
47A4xukqDgo89uqm5o7xMLbU6sSwCWmy1Yni9QwzAawaD2f12JWKiAeicLNKGkn568uBdwIafndI
n+Nv+XXiLMJ+JHk1TwbYgQqjC+CFgGJHdagnMWBxEc6CxJzLOCn5rFaP3oAuyQLJMS9eGeELQUW/
+yQqEp5GFOpNf9AVoFgxnLSMH0SN1UUgxSlR9JuB1Dkr6usK6QOFjV+PUK/2DHsk18V7tPvrQwYQ
Hx7jwQ+GEah5DAuuidx4b++j97Z7tVATAbWsQANrbYp/ADb8uXuei+R2t9lbtPBLXF8E+YZ26TmH
SYrwvo8/kOk5Q3PQ9Z+ti8oT2ge5D5y+TFu92VqNCtR/pDxeebaEltZUC3DfBl25pAs/7wDGDD4m
o1rt3Vgl1ZRUoYKTKQEg0mKO0d1ZQXNg/Cdd8FvZ54TjfWrUKbez/jLrkcLAvQuSZQfYRAsUgdbY
gxZlDiZhwgiK+ofdaAUyZ+QN6ngCpEqKn+b7WYfpZnpBuVEsrWSPMt612JcMLf35RObK5YG1GgpD
Mk3wkmQPQ5RDMr+eag/oRkKokJbRXW778vfvJE0Tz7vY7KyRXeKFs9hT73WR9KHD3YWEINh5mmaE
At+AxE45pgZGimmnlCk0dLuP+xeMl9S6vxeGdrnTGkJBTqPNpOQrjEqOz8PAQjF7lHcTSlIde14v
ngDirnYWm+wvxJKXuaAHgZa73077wGEJObVQOLHcyn2D5WZZl/HZs3sNzlrlMphVctYVZJh7fd51
4AaGqapY1dqLS+4szxuzVNzE6pViKysZyKWwu6z8jFzoHrQ/OvNXhKqlIIUFxH2Lj2klw3g+kX/l
pbLqRAqvyXDOHaUiZv+Zsj8NTkqfJKsKLE3i48AfQyxBvEQ6VixPjiUy8YX2wrF5MKXjzXBRfNmF
pkGadw+h8ppFHmjfN0mXLQmDD4NYtyShvDw6g7Ixx6hVlHKWNA/O1NMDSb+NiqVvZtuh3TJmKLip
MYUHmQcGmCBfD6SSk9nzYDp5UIq36ZxUNyXTopo+X9LAa5S08W047KYxOwPVe98O4fn0OW0fT3iN
sam/uGi19c5LRkO6lMc7udobCnnGr6GFk5olEdj7Es0G5EV2Q0ZsKQfQOC7v84Sa/UxRlExh/R5X
bVLteBaWuZH+bMudOLZ9Da6DqaCTdF9nNuS1j5oFz0Ldh5YqI5rFOtSPUGM/Ks2MFBoday0V8GCT
RgLM2VMn1PB5HJr9nWOsTeGSbR61fbW6KM7VskuZKE6PCvjnHgQi1JPYtr4/mMgtHCZhJwsNqAdZ
5RlD561r4HGfub7i3C6DbGOw57TeaSyFHvsD+gYGqxEAmLc78G1IEX7B2vK4VAutiyIsLYenjqS6
/7lIEo2cwzmKMdxNIgXuVvwBuUql4wE/zhl0qhE2nZl0tBr7068B09p1DU9lmVghHfGqAQiviEun
K76iVI/oO3wTnFhXW4BmCtT2iljKdx+phP0if6PuXUpu24B5zNBIX3OOTL0xyyPf7eEoC0ApzgZp
XBx6ci8nAKfFpkBBYfAAPb7y5qnzuxkOmpLHzq9HF/0/5IfQTGOZ7mzgUgPWufZVDDOms33hS9S5
MhPzwDhqo0suoFjGfzIkzpAxPIGGu7NJfqgVFD5ci2p7Vq5Lljh6tvHzse4JuIzYu3g+qb9eawmd
1wlfQqAlaZcC/YdTP3kRHkoeK+Xdzo2ZL0H/GZbTQ5/qpTa2qdcMwO3s+toBbUmJE6O+C8tgVLwA
jWAV5Oe7WZc4fIOuyvqFSByhtfHlRLZeq4y3RbTSdC9izuh++MBrE79wjtVvW6DJoaxp2CXp1dYt
jKneiKbpRHzmLypts/jx6eBmFx+KLh9Q8uJwiPkADF3KdV+LtOLZddqAkz682XVeWLgL99Fpkhld
CyBwjRjm0m+dS6rJeEX7RAsecWUjbXsouucWZgk9y9N5noHuHOYO2CwNcwu+XcL5h94XDkBdm1Yw
hRMn0gx9RAcHghcs+KcNwNhELfC1WForspHRnX/j4Txs+QTxHGouY/xoBzarO96zj+QGlyfcoTPg
7U+MdUgk0619d5egw2g9naHN0ATLHHN6MZSnBz9gENa0OcCAx5mjsGuIe1/l9lUK8pu/VpaPn0FT
yZ6AzMRNuuUv+svak1b4nhy+xJHMAzTuqnl+aiBKh9PCquZhp6RpP/Wh+3lnEpZEDEdM9G0wu1tH
cv0ZlttAUDFX2ZHXjEWhsPNdeADAfjTAVFhaU853LHOf+k9HzZ7Zrtk8hrRNN9qrfroPv1286Cf6
4gj3sPf15uoguPfFhxkyGwOXb9ps+Nc7BfW2LHIpa3QNGnfF6T7KaeE3QePsA8ZbD9kekMbnoGqe
re3wL6zBzobtGmDwhFNtUnv7IMg/EVlrGCNj/PpZjhPoX66Sju/HsqydyCVGcFxfIbREz5mTNYKr
zA5SRNqFeoWkdcZvEjtIK+msRN1OysjOuBCOl4n2Y/XMcs40rm+rQZq7bR8wowIKbtSZNxxFaiC0
t00iMTPBjJLrwCoyD0+jcFEDJLkgimzcG7tklF9im2gccPPrbu+49P8/kPp2M7Rr1dNUxTcdg78d
Jl5JP3bU8WAr6FqEOHYnf7ymYMx5XhFTKjLHHwjbzIWK/39gB2gVsMDhr1E++S6KtlyBsdwktErC
F8wHSfGNNDEEp/0YNynmFRkUgDOceoRn9BaxbwHXyNTzsSElT+LaN0/oVoDKGzVJLLVAUtuKHwoY
XpYmA0mvHiufHZVrRkWGWdP5HjSG8rO2ZH+CYuPCU9O+Qh2sE2dZYnPPmaJpyL20C1EdPM/b4C3C
AmxcfkLXaFVNWOQWtsZVCbNJdyQwkZCXpVhfkMjY5QxBcOCundNSbw3ISlZ6UjxT5yC+s+Jf2NBj
jiZp9CJx0ckqj5GOXREx3pufDMXX4NXPr6w/e+SADmJXMtomG5P21M/CkhrtpK7Yl1gKKrsvNvLt
Sv5WoDgULodMltJxwwRn0giecj7/3t7b/c+pjf5BW67zb4kOWGQ1VcfIXx1MNULz4yCVrRAt6rQC
tYQW3DMIT/qCvoYqYU0EihW2N0xGVVQ690/yqXq60zzZZaLOtE/bMaEt1c8scr13p2zLQU/ZZFe1
pSUa29ANpL7pJ/amYEz5Ni0gU15rnqZrwRqZetcj2uvC3i05EkeTTUj4QVub3+hfWqGYOE2CoHft
FlHFQoMEv3dYfQQuRNeU7SVHhTX+2SFoGu4x3UvwHFL+qzH41YHCGsg9uHJXnRCSG3G/Ws2fqI1+
cQS02bd/+tRLQM9sV3MhDVUZtRyn+Mq5SBcqSnPNVAdXiqbJnnxg+YBYQYlFZ/WeHvmKKNq1AYPH
STObYRPCrNZppugVMMeKnwzi1V6TImeHzZ+vtg5Cu2XtA8+PfgqBacHi/o0NqMLcusyYNt108L8h
mh8GXkbgozk2Tbo0wnx+rpeOQlgCsbQUijkJQVOlB1P1LnXmNCn4X+83Va2OHQfkEbj2Oq9Fa4VH
b21PxOE3TLzQCb9r7dS6vBXS5uPI3VKhppBCCpUIm2AJr3MRs0UGuWqATdXRb6uDCYsvLUrWKBlk
YYelyg/Dtu1K7RlLenBVz1H1iVSEbvLnqavM8+99Vto2Fv1T/tCmQXUwhKpT/vzhoRBgbjUEu3iS
RCzhIHI37dViZLpBagmvcipa4uAOi4hxaOeBXAGf0v9VxSzMiMYjgDJgHEDt7SMNf+OvIDknGGyr
3/Ryb8xk2fzYBLUbTop5Hzmt3y0nq38b+JfS9uu9C7fpcwb/LL9GYqEuKg26lu0e8wUno5PQR9O0
mWP4Axlaa1JROymC/MRzTPFFADY9pPxJs56uuN1JoS6OODrIUZZ0dIpLyFvRN4B6vbNmdF/QZhAd
3XO2vKF7bn+msU5btqyXNcV4ofBip8LSLntO1+JaHYkzqMMNOj3qTY3u/p3CnGn8d0J6678CZ/Za
kdBYOahWDRmlEfQO5ZkbzB5LHCi8xTofIIIkzMGQ1Z2yA9T8orTRMhDDDrb5WrGXM9aqYTyxdkEl
2xifSFY3IAbl4FUX1Q7q7CrKhUflCu2CzCPHlKhMklryjut7elPikzcd2SWiKzjE2MQwhfJQ0AMG
kGKF2CGCB2vSyU28p3f3zVA0CrjZjRz+WV25DKnWUH/jBiEEUCypxN3gr5SudCBQBHUxmlxaVes7
dZtw1Hs7edhpjhHYRqphTaQh3znhv9QZTl+4d+lLAND3Tq1tFCaYVhmukkbUgmPRqXxSWuiYxq2n
mOdXDL6yuJ7db6qswkTprkkLiJU2P3LAN+Nkuo7opNou0YNv/2BxSvK5l8v5OLfrrcqQj/BhBvoK
+Z6O7IBNu9vgzdfmMOyralzvFPCAEFyfU93NU81sibicmKoaWXbiCMcI8R2IY6kLHz1V/e8SooW6
OK5bGsnuHigeJPynGpVGYWmbU2JpnBm47K53CSjpSgLyCpbkKKVOC+jc4visdHAxoOxOipES8M+z
ku8wyC7F+ENebbzqvg7g/XmzvqWCm2aEvAhpAv1Lz9OqyKAb+fAu6ZAGaFH8jSLHudXKrEg34OKf
ykYBjPaYhRhcKx2ZVmlrNwqCeKd0U+I2FClMAq92wu2+magnyVMqouW5BIvsbXH/ktry8IcoY8oN
owgBmviPJCHY3ZzyP6iSsbanRR5srrtr2wngaYAwkCHFU282F3Y6Hre2oDrbn4TTbBMizGkBhO8z
gJN1sl88el5c9xgJKnFDuTbponx4Kvt7ivHOKRcx2dP5DXGlJDha0OH8AS5h8kcxf7FmtGSYGMvv
H3lPwKdivd3ATBFvJg/OjuObQPjWmJebgKrspCsZMR5t2n5MLns3jAWn5h6qHJqQH+Opl2ObGSmA
LwWhfLMOTAyaX094JYLgOMsNrziusfbPGciDU2w4LETM/SJr0zHHh4jr1DQC6fmlrSzLua3Y8xqz
wzTuFw/y/YnSFlnBRUO2KchBIAZkpGlA7v2SoCCMeu2fq4anqQvUK9qoGuiYBlPzzeQC+UMH3nqx
KPL/SGfCJWVEX/0PqettuZ+Bc7lr3tHSm8jz07+5dO0R0O1UJ8wBB14om1TMlGujQYNJNpQEujnV
FiG419ZJ1967Z94C0vbkRTeX5OVsfmJ6yDM0dDQ9s20l0+zHEAb2j5f4aswabhzc0ms1RcUbqIf7
4O+6CJiOhy5UopNK2N524jUVIalw6c9Zr9dt9l8SBIsICgdQMwt9Bdsa94gXQn3d+5AwnDV+5fQZ
WHvxaaHyV4LA/BNN11In0/q3yPdGGoekqGiIZ9xrGeWxPckw4snTW3c2d++sFvdbs8kNcBirHb1J
W8Qju/w4eVLd5G+BRWTgfmQTCl8yr5nN0qO1+2bqTIA0GgHpHTHF8lOcKw668P2c0n1TOhGOn/S4
kQJINge0x+Ksu6zGIwvJ+iyRqY8M5ISW9O40xOQbmJ08qUfxthtRBvSn0WgU1Qfp2uFzyuRoYnC8
vATp6x0G2b7IwM+m0Cim2n8SeC0Ny8t3ffIsaJdqtnvYyCIrMWP7ag9Ln5FHilyEEs72qz1ziiMa
IPRs4DWj7Fguv5mhfdJHIzMWR4VJoIbiqK4Vt5NDjYYMTxy21MEmP1RNVMJ5GQHO0A3hLpWSUICa
XGk1YEG4f/eJ7lJtQMUMmq1sfwFWYBNPtz7b2nT+Q22SxaK/ZsNjRQ2fBtGkws9ArQrpnzas1L+n
3whNyeoQ0Eb1yeNdvB4soiVqhBuekrfbJERYCYrGJVKG/iG8ICEgf88zbk9a5ePp0nciROniEdqi
ni3xLIOQQYgGi2IZTEw+rMKs71uh15on3CxJRqscj4keaVTE6MrSTYHHNrAwoDPdxQ482zQThsai
EUug4x4DN22jOXq+AI5vUj97FhHgNX6l1YdU1lLfdOAfRZT+F2ti1f2nXYVtSqdHzkoxsxG1W1IH
g5DxBue6Tghypoc70vGVFEL3CyspQxYSBn2DbEBBSUUGRhqXmYXZr/1FbL0k5W0tcxFvU35mhuOk
9KXF9D9gYk7a4bOwYCu68Qz4and7X7mS4ijS1sR3l6Fb4y0XA6rkV1H7fRmFxsBfWb0Tz8RgaoHJ
y6R+8H/iE4fwXvyI7msqu1PvOIiKUyW1iKOPuteq8+LP/PsDni8hjBp7ecipVCzbKQ7k9hMpbi+t
J0EhavHtHqDnDLkV6Jv+0FJMWhwrXvwpVMsdqPw067YITHDNUa+a9nt1dtVjZ461PefqPz7KGoJu
WCijKxYAy/C7TLkKg6nJrpGHuAfwGw2l1YDm5wty3yNYXAQ7kgqXZnqn7xHM0mdbjM0/mhM4jOf0
brZVhoFXqtenl9WBefBkdNw9DY3ANKr37xusZh3IpEGerGFU9AosRE+RvSNwJDSE5id3UjWzqErI
W2ZrKQ9nS0ckWKqGhlK4QnYy5X1CEwshFx+w/GZP5mxlm4F1qR5xTrMGLVEj01VeMw6eyTf0OhmO
Ipyg41nbCHcHRckSM8N6I37dz2jIf53uvW2EYCdeSg5npVZwNH0SoF7r7imipOp4aruPtkiSjQzl
lqENBs3Wez0d5LhXoyf8RK150Vod4a+mdHJznGLeh8XemFDvV0CW6GsRcXjZnGr8D5gY9Ed2K6c4
u4pLV5LcOUJQ/Z9J2/2zyXwDLmYvtNiD/ZQg2b49H5YOK6Qt1/OutL34O5U1BqieZAoZzzTFTpX/
xhJyVeMBP/7SW1khE+4LeAaUZU+8dyggBpLtkX2HmcaKVljxCuDiRmuwhq2r5lRdkvVG69dBJwcw
OWoYgovGwAUJ1e5byUwbhFpGjGX4e62BljSX6JKUp0pKbBfUpXEuEl77yNcvTSThxyzYkRtxDbMJ
AqD+hiNBjLZASfgftxfeWsNUMuKOPmiMY8Vuz20Ppi3HH0eha19PoagAzn9yL5RkGX5dmjMesxk0
Z2qrDk5HHe5ZrrnHjyR4smw8adlxg3coA0MvU7wnSGd0cHt7Ow0SfCISVKvQ0yAnXeHqExg/8spV
1KkE0QXvWL+kptfKwhLWBLIcJdx0bLl2a0a+EyPBpiut04Rg5mjLb2I7vEIj40OTcS8jXORrpi36
51YmMYO/8AV1mvy+Azlr0d9QFApmax+W1JxT5zgtTJiBSHSIk7bennkODqcfTKpvDgPklgWU3d8f
bK+rCx3rF7OeA24dGotLRa/RVCaliWjZcYzddrawf9zK4cdxmoRp5QqE87owNKvaYvWJeOxMDaWi
vfBMhvRFrGM8R2mzaZVT/KB3cKNv6H27391Eg9k2c6kdlAqj8bZrkgzqHPVtaQ7DdrIDe6aU6Vcz
39F17Uo9kSdYpm+9ijkuQHDYqpeu/v34fD3chO5iCia/BlGbogT16yOo9oYJTU8w6biZmMXsB8cu
aqfN4GuV8kJ6/0+xDwPbkZ7S9HUzs5gJgy4Iz7Gib38TglOY/3R/9jqt2XPgVRT8DUmp6e89fp1s
2Yc5BV8X7tfcC3s8OT5oGs/h7Brn5k5iEYsjtcgx/yCZBKVrgSg6yJEUazhJn8qvC+LsyAzbU9pC
YU7IMFvTIxH3CG26p+0OnOdivi2IG1WxweXYjVqaCN7pOfTGvzk74xQ8+TN31w1/5yT0wRFzZMEe
BgyISUL6BneY2TIgTNg3v/M9YI1COqNs/wX79d3sYk3z6/UmtDq/JSLjO3HFXotvcYWJ2wEmtqOU
F4Xu76/se26kwMTcLkIYNStpJFl3VyX+D3Ry5zhhPwanbmLaM28CVWCDKBUAQGYP/N9oLy3CaoDG
yc3EJ5yJDRELpJ2oWbCmn2pdTY9HazJkFBvCv+EyNVkNddcH4QrWDYE987ivL2J0VzC7oUH375CF
cprTUW6dI1e/P1l98MUNacSifiC90gNpSTOsSfLLh1wxtt3kbSB29/k/9C2Yq1/WO2TiZgEJK2Z7
AHYABTZg7ijXrf2kkbXqcUkqSUP6ubymEETEmViDR3wVee9KsLcIES6eFO9Az/sCn9v0kOMYWfTA
rkXOHecXwFaY+860YUm68D/fnrLjXUSomwwwLK0cnlnlGx3bfOzJ8bCQqpr48N+frYiQvX5zzN1s
V2QnqTk8FfxIm+/LiAvjc1O3BAVPe9AJUHbD5TMeXj3sc6lZ0W6gLfzachiI49cqY8x/s+khdNjt
nUHinNQrNX/26SWxUJkegeO2tVLd6xFAyoQ/oy3aclJiPRJbOjsPG09roNSvAmb2JnGHBrs1jpyM
zrJWKu1pGgMHimvjL5CK9k3vA6FmY1/XtPdAOfFsfERbYieb5aa3oNNmjEXCC3ZA3TcR1hoGkdDQ
Ou04sHzt2skaVA84vc26CSevG4doN/DZizfz6cIFNU6RMecRT7yiOLG4cfnsJFJzHaWfcDTidYDf
qMXjUG8+KuOxvLdK2tEe8HswgP6+RTNzJDuN6uNJLZzi80WPbrVlQJF6Zrq4QirJ41ISt91F2tIR
+6trOVPIEYPa0DLVsDQU+hezsc0JRzxTy8Zj32xskPWxvqTzAk4+04VJqQXk6z5yhI1LOWehAuuq
2QKn6AneZPLTg4wb7HPl71yI2BRFY/EVYvCp5nhkDldYwLsbfSG9p9FdT+8JfkdlsW8fa1fkdAWZ
7ZUrnHRm51Yhzw4hRluxXbVjlg3T0tLGrd+z5C/pa+uK4jxmL5YclZAy64Q24Z6FB0Cy6VnOBRL3
Gx+/IvhEJZpGUi0WnZnq97CRoXmz2FRu99jk9KKdCs7l+1TuyPPsTNK5hRkOmm9KaOO8d4HuAJHB
zwTHATdiJcoQh7Cen9AB8rKosXSWJ9lPOtElLQ/wOkrCTcvWABqlo9D6USMmxkLeVcTYmaDFQyyQ
o2xm9rLsNN7bCEItMn22v3HAUJTm226NV95SI6+6jwrMZ3lRcFJFNvEGqTLcfoFNrjTciwxgTdW/
qWa/O8T2KTsiWeBhGy41bi4mIg+4ss2Yxk/zi2BUHrs4RUE9NWriqk35seSQ4j+StMSdTBIRP2iF
ur4YscvIlp8F63saKQDShg5kzqUWOkfeFxYHy51uyVX76Ha3ih8b4VvW2ToQuVAQaNHvDzPG+wGA
P6iFQ7zFBAn5cj6KoiACkQmMvrOcb9MLtw52yQD/I5q1pzZmLKf1rwE/zeWkp06NbW7sL13yxqZ3
uUeJBBJ4PNaRbPWlNNdwzzUqbubAyfxkVJVYrDR+AgQY8BBTkjjKxsSAH+yOuygPyY/dieBNvKGe
IMajM5TD6hrCkAdUvxVcryvum93WoI4dSbf02gFnGAIGYKygjGQs1VG8kUeTUrD2fGBJIOgx5QpE
OXsXO8NTfiEns9H3k42CFcy/QXeYR614TtsbXjeAtuiCOcpb8nZejjeUSmpKxFjWLL6JJNncyeSa
vX47oQEr4lx/l3PR3pJBmzolGN8ZRmbFDrYPkTtIVDLU1lg9co0bxsxo14nu7lEEJb/OCT06cGA9
F2z13EqzqoJxbFX+2ojwMRW33A8TJZVjgAC6qMmX66/ayAPHpbLq9h1/esZaKZ7igOYabp0gcdFN
9D8Wx01mGGfRm0LjETD/1bt3Y4VBcQ/wKPNVG+XqJ8H2gI6mwlbACUR4OzNsRIwcvTGm6VzFFP4D
Pu5mrv8zFDLmXG1LYeSFf0rjJq9tG5fkBsR8jCbJ5J/oTUXThvvNg+haxDOXWCb2KDWQzvP0uyoE
+scH6PY3f6v+H2hjYD2iXNsNUexSWO9e5JCz7iBPnCRgLbZ19eF/v2GDLKDHQNMnJ9XVPO+KJP9g
FRjq1Pnx2fvkTv7Xkz1PNqQcMy/QHddHDQ+Vlx4RuVsq9lEx7wvQdK3U4q+Ux7alzfTgBPIrhBew
+II/YLzUvkIzJp8FW7jhDpXwZ2s5/ska9bCDUOaOrKAX+EqHnq69+ozXBDGuWMVzuo/N5/cE8BBV
zDaL0gbXSF+aNat4r9lsvDfasJiep/at9Do06TGw2qpGVDivA+VWsA0bN9+ImhO4nNioAJ7zVECB
uAWFo0m/nBasIevxlGyZQDFMLchip3JS5ZaW8MUWsNl8bwLGF1VuAA0PFia6+ZUxWxe5YY6bchSz
v/jnsubpFZcR/ip63mF6Soa+SLKxSERg+uFkMDgY8DO9Ihun3BMMHN5/neroeGN4elo8scO9mjq0
Tn5NZf438PFVCWWfaW9u1rqbX5FGcITqSPEstNZsaubc9IwW83Djxe4iKACXcpdB4Oe5AOjq50z4
SQtwqC7zgrvbfj9X+F5bhcmAqyUPTiiZEqnFyUe/sONa1l2O3z7HQz8BlMBKe6u9uTYVoqIFxt6k
tG+TeCGYyZodVJX40OvMY4WJAEG/IwJXaWXCFGPKVfOvtePd6hWGcISwl8xsxVeV0qcgWYVNLZc/
YHjiArPmiAHVWv3NY/ZfeUUZ2tXmf47XWa58Rd9wMpaKDcfx/HlvYaD4jWGm37INzByq1ClSuOjR
73zvI36+0OstZxkllVcWySSbfQmXNUyH/YIg8xr/w3ygxBZAjmKJMbAO8GmYZE1HWsnCj5oYyRJN
0T6fYO+T+c72AcjOdAUkCxxdALoKoEm3tGasBI3MLpIxLlmClFIBjL+FAzawTjFXEdVtZrNHr1e4
uzxx5Wcvdfz+kyqTwNsmRMtpyPTDyj8mG6ODrAD8O0e6n7jn07rRX0waMg39P+JBavBsAcdiW9tN
4iJp6Mr+o19bi0TBfO5VgRp3xw0NElAXmOVSIy++ZmhAeLPrAGmYAHi83AwaJFuW2FFa562lYDw2
5e85ZpeDYaKnd3SAyi38QAkMoufX0c3MaKKuvPLBgtlqnpcvjouUeOt6KmjQ1B5UQiLD+ip+YDoy
7MDmRBwuwq1pwABEAWoCGtU9ZHDW9CgPPRx5q9ghZfmJK5B1+gDsZCU+ZvziYMMVaCocfxUSwiv7
0tlnLdT5+wHzrdw5n5HN5A4AcUARjsyK9xM/p/k/u903/3WagvKdYb6P3ihp7k3d2WUQTG3XuxOF
sICVdvlSq9/0ped+J8Y1qnGvFc8y3XrIqpCnDdLkT7OLv/f8QrxQ8C8tcdk6MX1bP/LWiNf5wQV7
VMGlLZ5B8egLvgaMMr/+D2jGlICvPkInW7UZ2w4GraODAXaCoky2b9yMqo3RZvvcnB/CiDGXD2Z9
mmIRqy8Xcx6EuzkS8iHByTY9Gb1Od68LMu4ra3bv54eLR1+A1tyYYe7P3UJNmswVAS9LdH+fRgSs
iefSJplGw34+q5gk1d9Ug7KAuKx09/UbgDiT9MEjk704aqZVFa6em9Frhud5Rusbu6m5v33GrfsX
j/5UUKXARl+/ZFbvRXNcT8TKCillb5cKHes0qFmhWIS+9sD7fWyoQKP8XGk4hMUjdzcIYrzRA4qs
jQWCqWrse4Qrmct7jefjQySrbg3T7U7WnhzXoA4W/OXDkb5z7loD4zlvrCGF75vnTjdjayNR5hBO
LAe2aAjsNAEBC2QWGhg2Btad1aGA/e7K13Uk6GAS1LGtfwC9Ynl+pQtP4fimiDByV+TkXztzOGBS
LeDK8GqH23jWXY3i8M+JLYflfsmfPf2CjqHRyRSwHG/Ef4wqLrJnlmJb6K9ooDuLR3dBB0slAQNR
1+dby0vN9FP47FSAp+0DMJdkJWPEv3/uhp39XLGSYutoBi3XbPKfYdzz3ckEKd4a5MjcaeMhknyu
W+/z0D87WW97ORKIdeYR5cdbHzcpiAjzNMJDOsZzPqm5ta/RaddLgeUXpBg1CYUaMu8UYnvlrMSO
ZAym3lfRyh+ppF6b1JoSKbSBGJkHthExEMiyOf4isni3yLf28LEWZLREDOf8ZyI+UptSpKtaD/jZ
pgYFumNELnO+URUpda4B565CV9RzhZtAuCtA/H1bS48KRG5tAyf1mFs58vbpVzXXJ1W6G/JH44vc
zp4Grx5GuxxtG7/yKrCTGGmVA6i4Fb18Rnhg1sG/CyoaX4oB3Por8JyseBef83aGWxDshdu06Fzv
RkZD/ZlvgqRZMUFTrP7MXSXOJULO5JQH6m2rcI0SdYs/wWsf+2ENRuVFnH57EGWJgY2hL8COGqPP
9G0pfzkxO7fgX28BVSwh73Rt4Vk8j3NOza8hIx5m773OmOTjrxafhyy/s2LqqaS75YGggQd8uTfW
kZxqWziqHVaK0jfOHvHRQGc+dQRg7tHn+ViP9rodKoY/onWr9oyX3JtqcuIGbGLJlcEjDAFYG35u
IdfAi5MAhiI4quKrm3WNjeShsga/mXq3evsO4CcVzFNF7EpbMWIHyvmb3Ei7FlX5gt0yf5/cE1qH
YReqdKL5EZdWnhTb8uVZv8a/3TLUF5pliobs7bTQl2aXnSdebhqx59pV57DyxFDKsxoLwFm8Vx+G
/b3jEjISvk4puDv+NewQXhdQGWnkmrZEeyANDHslcfTG4kjsfB+tTPpmKBxhjf8BGYnv0+0SBxN3
2jqU5pjGPGwnIlRvIK/mue0eCU0+DljdJvJXnB1BlmAkIK0GCRJJDCe8G5a/LgSWRMHTVjRXOoA9
m+DGJ/heBPPMs+K/W2dm/dU8M2el+o1XWNbGkjesxSqXsBkOmbuI9e+3SscAQ75GUJgWMdwg3mtG
mH60aIMSv6E3C51lZhKKuig1G27eujQJquBTkOQjOiYR1YRwRzb58JNuttRHxWCu2Hdfz1zNaZJp
0gcNodYAtIKWKKdnyCndV7wg2Th2HY6B7agj9LPUZVPiAhFJsmKBF3dKmBxqWBj5snRE9L0pAo/x
D0mKPIcRjyCp33YeWj/hUzlTPCgBW+7qNycxHY0WDWI6bkMpkcG3aRDOoZxIUs3XKkLnj/4pseL/
h6r3+MSI1S01CCZaO1fdxH+yZPGnjb3YxnD6jg20GePklqV8m7PtdKeRkjyW+5KVhcgZTp7LK3pq
H3T4IOzpgJSq6Hef+P86PZVInL/yDcw1uc4t6A4dypabW0As7Jl2Qh0Bl1nckqmLkr6xJ+xac35+
HsUtuBzBns2Nm3ghShuoWCkNI6KNStutBHudZOOhj/kBfV02uKJlxWKr29GpGWk40JF7uQ1+8+RV
pn9sL9ULSd6ersDJQlw1F3VStQN6UDTJlKK0s3koiS5fMdj5/xPEZWSPHwxW8LAwEPFfLlRr6ZPs
SUTIhmLP/QLQ8pb0vRavmL3EKh5x1m4AgCpZJ4ORYXdqBnO8wNrhj/MMzh1MRRol1uPCEb9B2pmN
gIkj6Cmb4OE9Yll5hYc3DS36bjmrrjBRHmyRr/QkXPVCOgOHRgl2s5GkmSMc2U498dXrCDsxby3M
opMxmfBK9ISxvFOamhQmLyacaXfot3i9J0WVmO695vTgmjzvMIcHVHAvUeqNDmJoYd6qIpJGwH85
y8ZMj2Cz/AKGNaAT6EE4SGqINSW4jzlrxPU5g5w5qcw2puFARo0HHGx0nQKHMMEpG1vA6tXk8doR
SbRThpW2M2ryuMNeRJEsgY6DUeLeaF7Z4ezoSl/nN6pwngNWeWoHZLwk2+hudUY6l4L7FlYI7iOa
i7OH+MKcBkUteZMWw8PwkOpdxrkG/v1njO/ztN3Naob2K9i+mBpnWp9xwZ7a7UsARhkZk1KYgsg1
SLAVbVj3ldYMwlxD/j/el+/yiDOHXfLDmlhKA7PZwYCo2aCgfUJX0ozNgydx0vt1R4cGIYmw/qLp
36nSpcE4UGIWuSSfDG+78Mdf/59flljZbEKFSsHDaKcctWedbjqmzuxD1SgNgitxju+aMWpclVZD
21IRNNoxR7XYuSChS/egkg5YBy3bSTocVescgeAI3zJ5wHQv/+mTPf+ybxyfbGiPOxdjccRsMWHj
NYmXkYkLzsXakx7IcQaI5Q7lGKWDf2Y74eBsd7R1h9JXcP105Ab3RujAF26DWdyTV8SE8wUf27NS
krGNn7foFb/1ujGl8DV0MZ1XvL8ir1VGRVP6BEctiNQmk9w1KWgjk/If5sGzokroSD5uck4VOZtf
boiD9OZmf1eRaDtksddEsjUJUOhMZp8MebpM4f8VAcKapCzu8E6TnY0d+fYs4lciLsnIYhK+OKnx
i7WPCgwJI0lE6BSWakLp7k6Rx9hOr4vrQP/XB/DGHFX91eyPWy6IycoHrX2TssYLbbebcgu4ggFn
6WK1dm707G1bU5pk8tdd8xoisRhUNpEw7EDC0/mvocq1w8H/1DrhK5ftnvI6xXlxxZ9SScjkw0wS
UNvoqDHfAxuk6TOilEmkkZSiitlr072vqDC+ZGmbijH4h0joq8c9Xln6UOJxZGVwqEfDPwnEmoEz
U1etd51nwp9xSEJHS6FYROrPR2eAa+t5i3LV9qJQCtMvDIqc6ttwytL3430s9LYjowcXruIooYru
J301SrjoXM60FLrtvZa/5LBZ8S6eG/+Wwum0LKZ63hXSb6MTTACXOT/lEIHDDDAHNiFar/PHBmLR
JzJNsWISRES7hWLlCY/SMDUb6FmTRX+HsP4z1zlrwuK6HUXNY9EUrTrXESlVKEi/VKS3cLNd+LUd
08bRRurgpLvw8X3vZXI6l/YRky6P5FiehCby2SLqWD2gms1t7SrqEhgzvv7RvXpXWfkSCfsWHpx6
LoLV4kfLzPZ8QE0B+pZNowyMG/3b6RIY5rJl98Cv/WebJXN7VjCwaPfeea9zmyKELQoaV4Ej5axU
k0koTLLp/SRjRYz04ZdYrV31kO+gwfwVTUt6TMItDR3eRt8xQVHSj44fT2glhA9vBgnF9lUk+f7s
9j9NkZnqoA8l5JJAugPou/81sZb+VoyJapqrfsepXWxv208/Gbr8fe2PXl/bAnH1U6ib2n8B5hQd
HdG85kvAdZlI1MheNMaAltkhpygj3gU/WgK5/hSnM6rQPoJkoTcvwaoDu2gSE1olRG4v8WMQcGA/
edL8x1p2kc4xAQ/FYERS8t/WRb6PFxsbv3K1pe+Y+w9pFFf3CZS5LlELkBcd6zxxTnL4SmT182NC
zW5qQDSUdfcCIPNtRZrxXIaUpOEJAEmTfkyZFZmcPrCMUvREd17ZpFMUA/KDnL4KH7xkazaMmnDH
GDLLE/vMX6FynZopGZlQg2LgeOu7G5kkeg7ireOCfTR3Qf/Rt6jpRxpUdt3pjOvWF7/kLXHWjoWM
Hl6Gw3H2KlRFo7sFiCG8k5mHvoB/VcVJ/tTUiacQcaipIdgMsrQIEejN+t8nBcijL7GHhan0OY47
32BjF287uDYKhQub8fX69VWJkguDF7RP5te94lw3gRlfD4s+aW4P294WAHAwlfEBljsn6l1hr0iQ
24o3Ua8C2snVozUj75y/w6krjYA3aMQa6oiP2qK1JaTRU7fvfMjGFuOOa5EIz7y8XB9H77iQVixY
40jZOPaDwEROYjvVK41eJMBLX2ShiXEfU0aD5kA/CyWSDfs4G1nMy4I0JSKLbqjA/Abk+IscSpWn
FE/+jpE379kp7yDeP4UJPueGxexl6cUtVpQdCt4CGdjmToZ/9L5mqbKG4CFKu0fiAEZkiC7n5dXi
FLwNU8TVFK2Bj94EOTY2LRXqa4Z+ITy/byxjGhffIOM10aO4mhTMR+bSVC6YEzXeAVCVvtIthWq1
3C5vhZ0Tf30nP+CU8Aj2v0Bshjp4XnFqAmv5Uj5wzIv5eXmn3X2uWf9mB2DMS4np9vr0ZH2JdWaj
AWTncfA6BwRAZB/ha2PwmgJdZa+1OlrRGTpN7g16PTzV6ulI2chHx7W+ioUq1jXhli2G39W/A9MK
nFb//BNwIQQQsi45i9h/OebhvtZEnSz+ZNExxPU8Hx3ZYju0F1x+kvI0FGfFBiRUM25QgXZyqJTT
ADh9ARYK47VppyqJ7ii4QW68NkfyakxelRQj5PDlrzb88t3vbysUR/v6jxaZM/rgWOjPzubiar0c
THHZrdijNlBk/kQpO8+uX7r0/XmqyEJZc3/nPaEMHlHE4mMQmdG9wbaiK4CxbYczQGnlTqqXcsVz
u6NeSlrVjqIq+TDRDeFP+CnFe/rSwpOuK4NUb+ZR+4rOkfeWmtcmmzJdVlsgz/bcdigE0ZF7N+9b
ri9RYmPdAhEj7ShrQaFcdgNTRuiHpdFeQbQI9WpTh0YdP9a1X8m8upTSovEOq65Fht6aamhojUpP
7MBS+UsvQzj+LiV9Di4B5TMa3JAsWQrZ9kTyyhatyFap6XMm99bVHkkO5EKgJMEpOHdAjBZNKEZo
JhpCb/gfKG4eaIxEijj5HnHnW/l4BCEsbC1let+ThqfS64XTsCZMsQ6PvoGUHQgQ8qNY9NDdWfRi
r+6PAsdNFF6E1G6KnC6khOAu1rxoL4LlJmo8oW4BMgkm1x8F6vBAkTr73AgFEupOen7Q8bkL0h+9
saei+qHiWpKiWBvB8LMmsxpky5pOC20b8VAc+sFVAcpzWrUBwd3TP63kQKp1lAdVVwOS3LD4W+WW
IQWjY/FyL4K7bDTbhPqhT6ZFIxPiaZzltJF1urIdqA+ZacXREOeZ2j6+fyNZjvPwmIYJXa9GpZpI
0TDzqKMA9Jl6Xfu5GLi2FDu4m8MQFdTke2WYAdWyEPskd/CHmcS6QNJjWr/8hRxQwfS2GXNtryuY
LK4dsfL44droY8DJpEiG/CwsoXPHQ5voZxnShTgGmP9mVTZknV4391vqAAFYDMqhLau7S/stBVv7
F+oYm3stidA2segUnGMRFx9ERSHKsAZoq2J0w5J/NlJsSGY8weth/llWFSWlraYl1P/I7VxXIvq6
xZ3U5ZZjjJ3xWunkT56JuVq3RfECOHOcXkZ1foG/w0muARFDwSg5N6Y/EwTGBE/u+4hd4aKyJUtt
CSFnqmDalRF205Zyye7Zerj6iKak/7F5taxjuQxOrUqx7tjIYALOvbXI+Ge+0wNBBgLiiJfcaN6c
/E1wztRuKtQxEgSnciEy3fkfiHV33quBbkchOexMEL9SSiRrENxtGHkD9LGSB+QmB16jDtVFUYFE
q63Nicte721hQcmIoYHdSGWCLe1R8ehdV+QoUffVWyJktcMtj97EMLR1EwoNrOZhHqk/uez8cqBg
r7RjxMJUkYEQoXQHnazZfnouiQpUJYmyburGxqscYafnCUZ2WFdrQclxlpJvn8La5OgQdAcBb4tz
A1DdCzN3Kpj4IoAlM3bXi5LG274dNnqmB/k+2q8l+Z/iG1Kh0tNE77J6UdOBX7mQ6SUfdy+6X6lA
Tfbc/5viDSFvELtBG+kpKaU/7eL6khk6dzweThv+7v2tXVOKlTZyR1Bph4jpi4mkD64F1kwBNeJd
uJnqFL+a5Wze6y3OKAtJJ85Yj17UNzlxLmkxjdRctzx8fknlquwjuKN1CEmptG48yDXOh5nN2Tc6
5koIet2YlqtmilZ4ILbyaV8dp4XzJYSfth77jfdI0Qni1ODRzI/mptby4XUWuqsLiKpv/HoVYeO9
XdOE+vuA2x+Ll/uDs9V0ra9PiwvQR4vWnMfXW1KqmuKyKqtEumWaZjoiwxCi/WLMrdgifIwGkOKw
JcNy1cm4DATMsEXkqeOd84C6jfcKEdXRpOQk/eXbm+3VeYc9cH/cF/NRS8e5ZQUNZwCq5OpMkWYd
DOpBWUTA/zeyy2PWyXVP75u5mXisXpK8OdOR6lay/hnZhCFFtfAQ/7FbuHZ+oDZ+iL9goYqoC9Mc
Q2lfrHyOEUJj0Jq5JvkCdfgSTDNdgmQgFQbCpopQ2E/GMPA3EeSCANCXpxH+2kmtH4C48tTvxIB6
Yo+wijh3Yp7dcEc3G2Pu6cOn3DtR+t6TqFBwM8QHllp/VYK0ikXN6qw0ReEhrBwK3cL4F+Q2K2Y/
c85A0lHhB0PHrm59Z1gl8MSxeDV2dn3t/iFob3ubpGg9ySE6uBvT/+8CT4LsbRIQF6GkUxFqLdMB
MQMPr/0r+A3rrRF3Op6fp00kr6Sef/jW2VpVmi+HYQ/iJTRrlVdPWe5N7Cm0bPaSOu8fl+nFLeFy
rE2CQE3hgsmV7R7BP6Gsc4Me0DwiFdm4N3FT1WQr8QAhkZI2P2ywUFsR5bbZu33EWQ7R7wf6R/2B
EvGRWEzNVKdA3FfKI4QId60ZOuoQC8b+na35fX6jRHLoLeFnzDG5vmPhnNf+Lqh4B03PxE36eh7s
P2NGpPQKGzUG1VBLeQ0AL1QOFAZyOiH4FHgvDNrQ8Y5CkUUK1gBbaEhNM3w2Zq8sNjdnpNawZc/2
4Up4PBeLuxfsjalclWUc1QLCHFJe7+6cktq9Gv5TaoPU0v9J140Ng/8rIiFRKkyDsLO26+Ff/awV
NmKFZXqq8TeezWpgpEQymRne5+p/SYlAPiCYz693t2yzYaw3sFTYoiA9MYY9oGVblT+oe9JGaCWv
hdRdlOoQvjm23eOhQ1oqcUNNaoUecaCDAZDcWPYMluiNrDV1it15JnRVPtJMyEsD3/0s+3U+9Gyw
oJirp2Ze/bR0WnGn1gf0HHrIAzEYwHPUmF76EyS6DUo3uFygKNFYaoGrIiZj18cWuiu7ptrF6Z4u
+KMAwuj12z0hxI3syLJcsVmmN5NMhB2VFWfFlAJuD66MbD0/rttkoHlZx38Pp27vAOV2brisR+Zy
a9mrnbhMpyj6pYhH11AldR+4D/UCwy3L3T0vFvyncEvOV8IhTTAlbGeqI5un7AZbwqPnn1L/mu7P
X+k8vQfhaznLSj0V75Xk30ennunm7cTyUaQPUDn8kZq/XBXTfmhnjoEXDXU8mZC+ZRyInF274PO5
Y6AGraYgWy0OD4BN5KzgFzaGZ7HAEH+uqrZ5AGHSmoD3GGIoPf9RJ4W+8l8F5u1lpMcu6xAKE9AH
NbZpfv8YeFJ6+Sl7b5jiMY8Tus4zOrYfMwCU7Yi4AyXG0Ydm0pFnn8CJ+x/mgq2QoqQNjc7qJH/S
SLgo6suABy8BxrUoPk9J4eOguawndo6D+y8LPMM1vizFhaBhRtfSth43wTPnRXNPtl/JBbP/lspg
67JkeD8aj6ElgLA2TJhPeb/su/A/2svBK19DbecY8U4Ts7gWdpwblLl/hbks4IU+AaiEm2ZELOJo
K3PowrEA3y2agw6Zrrn+8P6jsWJiVZyf+HKb7V5OzLJLKzUq3PNm4XhTlNjeBXiPQyKPvZpWfWRa
Ix4d8KYrKM/gCrWZxdxmB+5+VzfcsrEPlfqHwEA28YXrwkBBXJTLgTa0vHrLgZor7DJaa1SYXK8C
yBDaHhb7QM8mfwWCMUuQhhf90GrCZImbjXntBp/KnnggsClNXQyvs4Yvpy6BNtEyAtn8V/zbPttC
Gj0OvGqpcVIrYU0cxHsaLOjexjDs7gvGQMIQ96LHYW5VXCSg3NnpuPg4gXWAxdytZCVHjGnhOPRt
ftLNaeqY7hsuHGKUVEPDh63zV6mQMX/vq30NQzazp+AIUK3G04pT+DcqnPoqqRqwnaDvEEFvZcRb
7FUhtO0HW+PxbT2H9remmks59B+pybm2N3lQ7OEK0cFanuKOA9ILJqWMDq7y9HUnmEJPhWjDX8Ty
YkOwxbX0OqllwNaMUcctS+egg5xrxGjvl2j7epjrsA6/mAW5iWNjMffjBkjRvDGx6LnTrynb2mut
cGenTqjQhaSAuiRIXwZ1g0LIuehcHdJ7nktlMWwC0Y5XohOL2MX9daSsSZvywRkY/drUhokWNPbM
r5oxsTxwXcYrlJ44HMjegTjzgiPu8dU9ysKKoJvkL3Nc7MHrZd8qjA+TKbc6+xHv6YfPcfI15qsO
Ajf4TeIcdQK5Z8KJexTcV/JiwWN7K/hhOTc6UVmng91eyumdRpCxf5Y4jTBfxqIuxmuz1IMJwHPH
3Gi+CKbui8qcGqLelXZSwCy9vULBgsWcqKErgAfMfW0VWGWoIbajbdVFMYVA7Fh4ur/6Ev/jW2Lv
X7UyVyL0/HkoBREajTK7CtaPyn75aApaNqQ0bkiTnzvkwNoMLpN63yNPf0GHkPvgvOrVO+dl8kB8
32M3yqkd6LGQ0FvbxAsoNDy5G+sh+nMXhlbiK7AfCUbDiPoqHTIqViC9jTqmz8RcW1aD5kp47aX3
KzgA9zWHcWxBpfnELI7lvAdnCYXTSyISjIKLTR5MiTTUc/0/EaSmzcsvEBT1bCvWdVyE05ZtUiLn
vqaA0t6lPQiDKBUu1PDx2KGboTrVzKI4KUeaCH5vF2hU5T125TlnOi+R2ddOvvi6C3YqBddWVcoB
QkSZxgy+wZE7zZqPPpqoFIINQyxccxy4u5yHWLnW9P15OOJAAkBbKwon7I7qo3xPPU9LtDLatHVN
+3hbZC6bG66n9ickd6Gd9OANMinr38xIXg3j7VScDvxFq7o4ZCZPVR++fqtGcqB2Dw+aPPXBzjxN
s4YJBCEhIY8yNwjCvvtrnBnCCRZaz9GNKipFUH0szEZlS412ZQ+Es2ESB9++SeM4aqS8jmq6hJJl
FQlxn/jnjxRBcg/JswzXe5fL8tVdjUbW/ysJzMVuULM6lFDYl+EsMhaB5XtSvY+c4FFVUyZQIVpX
HeeXWxMQhVGNNlyA5r7jrQYNBagw4SsxA25RGMuIIb7RO7w9sZhp9XU0An0PfvQjSMjHRwanwicb
8y/Ke8Ui9yloR6kncB41EFbYLhjPWQnn7JeUybM8dvgwkp4kJvJ/NSdtZyNQsLNWWGVHKW1vRRqm
+P7d5Qfwk8W7/NXZV0BEBT2MtwMOxtqn/heNFJq8G8YsY+vD3XBUqSZhNCUCbS6Ri/wRLlb2nV9l
l+RcpnK3UDjAgl5HgkCARJafv8V7gkS/ZsPWvBMcgnMhw/BAe7iOaeNHt2wOIUP4fzIRRVzsvFv4
4DUlFhBcdylfa21CiDKbBqZ0Ib7RgKgbdtKhKVQnqudIB/CoDNFvLkMCVlVMcz3MpwANGFJm8RlZ
iR8TDNx7AfhHFIuHXd3beI/zdffF5nzB9IQ/lE1W+NHrEDtGKpap9wrVRxNvLA/38wdLPHnQVFfz
RdEB4f+XCMVa9lIVfEf6YbNS1/7OyG2WvmPuAeTgGofLRjxq1ZixnuNdiRtoWDxWczi62TL/Ev9K
1IjVvcM0yce/16n2fy1yjD1a8gL1RR82LsIUh0RAz0jofmmx+zZJQ4L7ugwfxPcZOpSaX4LTHGqV
hQAqBJpc+KIz2oEGnvyrMJreHvKQvTpPN04rzwYUvMp9jB7j7HK2rNbc5HX29YXrlxWmswCYytZP
tUOJVsWAQo3jdW5x+xHsKtNXswnYROWcU6ksBVBwg3i6RHdgtpjDlHMPnCk4x0B9/+BLNqcT1fm7
RyT/vCwtolfSD548MoUZfGond8aj8Q+oF/O/p7XikENnq4yrjWuiwgCHTfFkEyIvmdY6tN0/wuM3
X8fnDET3HFJ6BbWFwZP3ZKMHNZYaCnQaxMAk4uhlDQxOfhagLtZj7s19AHwmosJ8YgG24Unn2mq1
sEDsdaARISUpmHQPKXNbrXUV1viGaWb3R3kwL0+md35DKgR52SersY6WA37zhGY98v8YiMa3IZHW
y2N1Wum6IumB1Uu/QX5fmRzIL1oJyPuqnvMrOtepfAXf7k/6IrJTmfJIO2Jhb13iTz2+dWkYAs9V
74I/NqxwBLckqftRL+OvO24lEVW06J+8wk0HGSoM2j1PL55BNO65NiQVRPbWJX+lT8BKdmBzF8HL
2e4fYLJmW/zzX3JOfFO6lIiohQomGToXk3EPQhxvRsYveYahYV+0qEoRtmsGHu+n3zywTWI7BRHN
CJCHSRm61FwIJNjgJ7DRwgS4QC+sE3rU3x8kXNxC0U3CI1S4nGo4u6t/BwrP/362U5ra6zjAf1Gp
IPGvtVpa/4ZguoE76qmF7lwuIuij+fqiM3f5K71pjMrzvYtQaZbNPM/VFxFmE7mwkBPbHtXWA7Bt
6p9e0G8cYLP/j2iruB5LpIbEgTQ0dnk39J9Jo2VrLAsZLaHiIHu1WbCbqDIGWZFOYMr0jkDhgxif
HVdqiWbmHgWxf7c4P2pSWN7TRRPl/Zvve5ll7PYMC+20fdnPo7ZXk+qQ3xeTAO5A4nzJGFmT67/j
x4hsRJb4HVPa+wogRdr+uG8ndSk9ZeaEuIpQg0CzsCbIZBpuZxzHcua1ny9xRzggGs5YJuzqVFc4
K62jJiczNv5YjyNFiAHctDYjr2ap/I5p3gFfTKAVWAu/vqppA52ovFRuCDmv9lhci8Zynsj3IuwS
o3BLfvgLoA6AidymTGNIvFZERccVqN7GkeH1Oo8Q2z//lbhrSyUXifosTuv4YdXna7HdLSl1iO3v
vZ5OOwbi0SSnzONyN32SHuRkcanQN2NwJIaztgWEZXbJyIZUnqq1NfGH72Dapepkbtnpc4eJYw0p
iySVy+350dbq3kwbPoRcSA7HV3F8K5uDF7b71dC2MYA9re3qob5NN2l73eNF6unMhH7e5amXDF9E
6sr7edSYmO3P3BI7BYJnN7tVNPzukjNpNCA390iQ7FXqapZipOYQZGyalkFwg2ARKlkPnWmC4JDC
k/ntPlteQPp7430XCQ/NA9OtLg4HSFCltqztxyy9/wG9Ef+Xu7+Hy8kNlSk9Gj3Jo7Thvqf0rdS2
QtbvvLT9sLFgEbt1PGel+CoHYvIaWawQPTfPMmE40rhabh9QZXc2rHmkaJJf42+IXX7SKuPghfcV
DKWQBUcslDypsk3uMbAtj8Bu0/KmzHnbzD9fnGCmz90ghp+WnRMfwPdzwCt/KJvoPYkJGAh12/yB
okJ7Apx9pBDw1m8N8EgRlIQfRXO64qRWhEZDpsnWtJsQJgh3HPnM8q9qXRW1E8+mil64a/FsRya/
wBAwhIZSGzM3Lve9ZntwGarbmXVWdBx6wI56h/crj0sVq+wzMW1rqGbvWFqFpFUzoOAqaXd00FtM
4FeItVJ7mERugdENVkCPMSJOvV367bFMY+bp3mM05rQaD3dqwuInL6rQu1y3X6PC3IVJH1VgAyMM
jHqRXCU538dkbRWXmgHQXDHhiDyJP373uWqlsKWvgL38dUoLU8ZwnywFoKohFbaUjq5DG+ZXTvv9
GyDxIDJLl/LWy7AY6Fx5HFB2+0+2GrhA2xb/4TeHFbFCiJW7PHePfN+GM+uSU4a4NC4l74cFOITw
rAOP/1Deu6RlvWs+GHvELq2N/WdxKnkHUl5Seokplj52kEseKRfz7TNVBXyecmA8fLiVmYvnptRV
i82uxdNi9Ox7976rnbXW0/A4yDRntoNnUXXP/OB8/Rgxe5sHqW1GPGSzmcLiXI6eMvDAW48oJ0X6
Fzit0b4p8yzBhggRWN3aIEDaZc5S/CL6CDgpk5ASOrRaH6DcR5KmfYx5u5NImXH+C7gS/xIkZcAS
XpnZY2U1rQkmX8h0hhmwxW/z7r2ULnmxVPx26rUjTerKmKVe9+HYRi3aYsKOtsbcJjHeAx1LEfZL
RVPEpy78luvz54305PEVYLuVATD2jHH7IKZGwWwv610qkc5H2wTWWGNTiitIxzEQ61fkKNwv6hdq
CZI3louLxlfNsqlcNzR6HI6cwf3Jp4c6WzavemaJdp5qdb2d5SypaDoKDsPT1If8h328HtlgxFRW
yuILyrk/FIiiylAC3Z6CcimiqScpeW1iPTdzwAcwVoo28kKiDtd3C+6ZhdI+pAZvA82IyHI4pnsv
BRkir78uTMmwNLtknoR7ej2m/KADh56qj72/OTiHCsZbjOrZwntB+SA1zRe1BE95SWLqgsM8Uipc
ovItfNRpy8oYTIF76l8KpRfJaLWDvnHsqFrML0Ajrflb7ippuBQHraU6C3oXFPlqRT1pfpOVuNLm
IvPFWJ0IXwiwma5XVnoYTn2T7DuYGVVCQUccF9V8EMj3rANATc+pv8Zc6J0Z9dpm+p6cY20hM+AM
FztxOhBMzK7eZ11YnjRdyhRHlu1m4DzNgofJxouFd7cZqHmUOSs5zPrSVquYvRuDGObV6YuAuU+j
UbLYaHBo+S8oBEJVwevaRNk/QjWHLDpwK9PSGQmNoHIZYG9jtSPzWOJoQLYI2d8sNiC/f7QEz/jJ
hmprSWZyQ1Kgvdckgig3S4E1WYKZxmNas+VOH7LOGod+ZxVJY6qqODG+xgrBp/f2eAYHQakH3oBW
AfRnbJcG6LEvCz6bjU1FQaBXbw9IClNjVL4mn3rUVpF8OkVkpUitE955QJjd5hao5UhM6kE2VKbr
p9vhKx9CriMIlkskThHzT2+YcFJxNHQKwQCMHWhuksgGZf5aHI1BpTu76Pog2cZjLKbSFHusnHOi
zJWDzTO8fAU/NSJNtdmsQROADYLl+cq5gMh+6N8knf7Jc1JEgLu3WAGsi9w2dcWtBQpSVKTvp/2R
c2lCR0rMH5hGBOaDSQCtNt+1pqXVTKIa3EUTgx2i0wzN1a6EpqJSjw1yZZzQ6W8WR3sUo+q8wJkX
9SMsY2ekU5plgxnymb4lc/R0BXkCNm3up7AauziyqT+mFLwWHVgr9RX8MusobvoBMd9jqVrdKQZD
B3SJSB2vOsuPjq3TZYC0o82bA0KBhaPE+eDiC36MI0dSCmby3cVUfbiRpUAazh+gTuG4pKDbRkzF
aQevsp1dlWYoxnRWXVoZ9Nbp5iNDnIvdYVBb5B6uymzUGLjMixUBUgJdrH+05kAOeYA02sSlg3HH
zw28W5M5tWfKGx+X87iy6fLTYReQAgJYAwKktu6vpJ2TwtpwudlISgl5UnOH3icZtaXmqkcIj8ul
FjE9Uuzp3w+l/itdhKqeg2hYQ/k+9xiooKB0mu2mbPT8AplkzjJB3dP5yr9ngCea3W/j7Nr56GJ7
isd+/i7ff6SQc/bC0RDOmxKtIeiDnITXumIjeJGXRpLLXYX/UDgRrvMpNU/SUPM8+m3c1RmaqvfT
yFQH873Q4aUujfnHHR7XkEqlgTZmQXSrXE6w3Ab92UQ3wmId70Ep9vz6M0n066IHKbPTMOay2CuX
trhN/Tl7fUAC65WPXtNgw6RtMGxSdaRVvLJT7HgWF5w37F/qW4wl/5FC8TJsd6qYcV1U8UYC6FWT
BAg3rRQowClmQxiOaYHWXujIt6UmJJeW1WC0VUSSLc2i9wxeyISw8M/bD3UexlrgDrXL8nJxHxmN
1/OfD9yl9oFrgjKk1PdQe5zcViT8iDv2K+wfywB2r1NMQK1QhKkD+DafPZkVo6zfwwaOG+tk1BUL
TBZTdCxgS8DgLMb8AVw2skEhHP/C3P0Eqt48vl4Tva7GQ4R2YIHyCNQpyFyPue6GPYxE1KVnvWKu
sFq0dKcuyGtkqXeIF9ufW94SzN909Kem4dXJfOdfUf0h6O23pkP+1uef4YbMq6j4EvcnpG8fueaY
XejywycIe5n+7lMSd/eTqQWZ7xu0rxdJYEtadOOt3GOLAE9T7tnwblpJ0J2r+DRhyjxqY4UdkZpM
xUmVrlg1upmafs6BuG8G7x30HHwW2fo19kf8vGmKwan6Yv+9dT6Pr87z0n/2B2SgHdXLxZcu80jg
u0RN/9yT7DxcNqTjoLYAwvzd9iwyqvjy4eoAyGPAr+1qoX7q/i9cbatjzCNXTJJzDxWOkUJtI3rw
6JdlEcBTJ1ZSRZjumMhYPO/rQpjD6txJ0lVxo6t9exgT78A7PI4It/6Fgx1oUUeHeRNlpShIywsO
T3T4EyWOUBwRZ6z90n8AkPjdkiYeTTGI87cinDLJWzs/eozWc0BNeSWTxDMLvTv3wgN4LJQJBIKK
zzQLvVVNVvBoHPeY8CDAfIo3Vs0bnmIESJmmyzOM/jzxM79gpbGE8sj05LGdt5antvXsW4Ci1Ex2
9crcm4M1A0OPInZ3Ih+SKr69FR8Qv3xbva7ggpUWBMUEraNOanhCgGXSXXVp7wUpKPIktGLM/ghD
1rlkr2dCuZAiMmL546S4QP+rgowx6o8+eG1eLQUgbeBOk6MtQsEFAfrGoe75swXY1+HpqnkBBJqM
H9JHjjeY1WC7uFEJGzYJyGv4Bn3cXl07BnVC5XwJUn1hj7QNqjJRSODQPKHHAejnXep1gaAJnDwY
PKpdOmtv9ifOWolFekrXY6tHucd8ZwD9fNmKPdjPM/6BtehBHSnYJPvWCap0v8FzGIuccQvlzyXX
a7qd0AZ40ON9dLc24As84h71pXz0zg//DEQKpWBUKfbTaS3xZ9kk59A6jCfWjUbUkr8BPZmDjEBA
nXRvlGEz2rAPnRlqPy1nwpFvJMiC/5PS0/GNiN6VwU30wVm+4sCliUgocoj0touETVBer16/u3Dj
DDm/2ycLJiRBKunMM8KIJEgHWCMu/q00qXS0vPsW7AghuF1IwcIwaCbf6hd9o1jIJawERnzphCIi
ZcZx38mvD50+DsP5krAES7C9XHdMs+oYo6JfLCV7EU2YhAaE6GiksKC24IqXH6cit4tsfoxOME9q
1S8faYiKr0qjnIyxch353XWwQRFJfJTvxe1wdGxM108/mVp1e/P5yrbE2bh5StQRSF74ZFRixuvm
MksTKiadTnLSd71x+h3mfEbcmx8IvXyEonZii34Mje9BlotOy1xx5yfOChPYIyVD5jsBnqtUu60K
xv/CfoFFKEYKnYy2u3ZOaCpGyWk+1SooeCVk+rCR8IM4K+YT2mNjM3GLRHIAimQs9iOf494Sgna1
6FdtVXMxODVy+mMyaSze6vNTOZQ4h1rESeLaixRH2CETf9EF/lMQ8dX6rwF7iGCRxXU7qTvqn+ZV
HIpgXdlotuRAwEHRpdazzngYpMMmR/eItch/vvYljSbAY7m8W1nutvWRGtsaDAVEziUZiDBQYl5s
e++27x01mbSxYyjvlI9CvzPFG+Emohb01c2p5F7etZ2/j74OAR0jOPJ6hS31DX2p9xXs5JtGz3Ok
9rh+pOO5/EvY07C9UV3lOlSVt18av3BnK6hoe4RHYFnFCM1AwIoj8kODRCyqmBMgpVlvuzEogOkZ
OB1GrstjqjS1LOLVE2zEzLq08BMNDEaLqKQzbHSVet220NxbOkfokhKH3h6DsZ6tUjH8LKu5Vh4m
B/KBKhzgfPV+P7O/7qambJay65HHpVFmlAhcRJzW8FDGf9xykbrzgK0LDB1niinJmRbUtJPh2oRA
W+4aEQF5qGdlVhP0MI7nfWMarv2DAV6bsRj/ZPEQaL+bD2yW+vN+IyAchyqOlz5sliX3KHqCRWrL
bCcPjFDfV9VcM5dTMBO0RcRXVw8AQ57HQcv5fH8lPhoYsJYstB7pgLkpgQ+4/2YKVvC2kxiaiDCN
BDoH1vYRPLeWrv0RotBG/ETbsAx1+oEm763I+n8eycUxkB4poLw68BPbGifAwUnzlgwX/PWSEUYy
yaXSqbcq+ovmqG1UYYJHysENes9xnk/HyVCejMrlXVJt96io+Tnt+UA3dGuWsU1w2m5NFaUjwmMH
ZznKLHy+E2d8+sayII4NeZM1Ie02knIVLcv1TzUYj0a3v1F0aSL7LPCB51V/oTi9EdUWutGi+gAm
DCKoFaZO7O1KJlJz1J5341XbwYHHVtjQTqPPVO6v43Hcb+EAovfLoy/o/AVG8LzF4OltCAk1TAW7
AWq+PGtFN6IH27uxFe1eXwK3XV/h+m6WiKyKdj9ylZsrUd0ijOhof+xq/BJtKLVi+nXzCKtFkkKF
r6dMq/tPqLWd/XQemSM8pcRE/ArRi1I07k9Iafbnp7CreDpF2hWWEF5QEhUf86kj//cHix0KzrSA
TX0ArCYGtsm6i21N/AwIzvT1v7MYCURIKHpvNBuJBCcM0+NHA0yNx8VyB8Pbr+1oUdg4vet+vUGI
5CR5EyEXkE2iTtEK/9eFAoDfOrTNVUe4YRsSu+xjKfFnimyd8kw1C4/PtOG+3MJZAbj+ySbN/RI8
wZYJWWSimKcTCPAvAFHVeoguVvWsThLwldAX4ZUhrTye3jjPAVEaK+Gt7mkVTXvSKLPQpT0WGNNj
ZfT6LINaXGYCq8ogA4ns+VCvA2VYtHBz7Ee/8ThdvE6oOGKE3zC4x0fjvF5BhL/I20COTgwKGorF
XmXR5CFKuP9CeJh/ejiEPF4gfjoEAaAocMU9qQmIqWYkscGHHmIfKODZtrjgN8/fAOBxGYtstpMM
Wpcfn75dpyD1SAJuR+FzkJmDJ0E2mgaLGOyZoOXJli8OwnADYQVdCDFpG4nObon78rjeJTEw6dNQ
qQF9HL9djxFmZJwVtFL8loQyF0tRYwTFCK+IY1ZR7pwAjtL6DpTlZwWar/9z2QQ5WEo56YnzJCIm
GaMGgQpitXmI3jmbo+C626NMcQYG33ob+quHsrDzujri8mYECKt598nZcnDH2Uqp04p62YT6jf7P
AmfhWvoxXGPYPmhtM/XCS5ZQJWETtDnfh3I9/SD9Dr0UwNjICs3lEzLV6cSodCP09vj2mZ2CNF+5
ttwys3A2hf5HpF1uFIKCrmoRlcLVEHFEYZn24/Z0Lr7/JTBXrf16AoOiQ/9K0/VwEtG/sx9TD/vZ
4Wj/YCxE2VSqM028N84fudpGFkYGSGJO8ZdDbeyEeDEFxAoYpDcZ2RsgvT2oPCuxxC4QF9sTZAyk
OjtAWAo+NkcikeENG4RL1bfnbjoXZSzK0FOi1ELCqHlLT1/RsyikDLLRMzfjjLfdsexc+fHAlsqi
EhbWhzuDnCgeVpRsbN8Scs2C96dcLz3Xyb5MhOA963WbkFV9PzaeLUz9fQdj++2H3J+uzQqNgdVR
amgxH/Is8OmXEd4scY10hnZZ3m1nk1zMkAS4haxE0+t4aAIlwVv9N2hsYuGZr+vEY1EOIxNr1o1c
bDMcWimzlWSLi0XjkwhYmtIZ05sfVipZlYWV6kpS2XHf/2VLrmcNz1bppkrXQNMf4sebdVjBakGA
jyPsIEcXfVmKdDK0KC1+g4kbkiHljrlKBkxSPPac48vc5bcHWm8RkKKEJ9LNDQVAK/F6nMXETdQk
H0P8qJXc92MQF7L92vz4KW9cO1XV6CYir6+oMAL18cQzgy/aEKAyo4l8sPt4Z+XsCR/pUs+TI/Q5
esTGdI5nWDXwYSF4/3d7UfBytK2SDYof0OoRsOewB3ZxQCooJJVazmisyMDlSUOAYWp+o4eg13A8
IJAgo0ojQV7dSv8qDZh/m3uu7Chnl4T6IgxjvirJe7EM1z1mR4GwLXiEzJN48d1ye6DjfNI3wnFX
jWinImNcYbEMOKaNO9gi8Tb6WTBjoZSVYtGIG7vdiHq5rxSTIna8jw4cL/1oxn6JvW1RcUwJhQGr
vSITWq0thkxi1iidnZd0BSh2lunS2Ya+KzTQ7pdCIdFWhqY09mZA//WRh+OGoeOA48v+21AHatct
vE6aR2f814q5ynsapj/yPVnyis9OCL8dl+gWaeSUpUcn+LxKGc/9O+RVMbbAhEkx/FhEABOtjU2n
GzKqrk9MdvXZjxJYK37uxJhQegApV1Spt3t6dQxneDuw7UPUjoH2CQq1OT5tlbQXkC0de9G4Eqgt
pQGX4hNxCYHScTCh2XIAIuGTwTLMjKOEj5edHm5sMcmBHqyQ8c5lMoshI2jSvrkFhWR8Cd663Lqm
FbbEvGrkKcPSmDpKR1fu80DbEqwN4DaIT7nZUjiQE7rFhOrtCtISFtOq/quyijeMgPgosaP1LKT4
5eF0wjCXXVe24mO055Ckx3UGgdXamT1WyCQg11gTNefXfRjQSi9QKEO/tc2/Fn/zoHedXHHnfgmf
Eavl1QTwXNJWCg7f2bvjPLEdOGBf+vCJ1ZHzHt0eH77CdsXHLFjNMOL5a9LqW0I1b6NyoYCmojxq
nrQxaxymhHjzkuumjpCc0Ky4Ivj5GUgIg3wARIr7G9n2agzNwUa1Np9NaTwRfczDj2Uv5aqs++Df
Q99CDAddR2GHBRyHmVedVZ7dPFfNFcgq+iUE51c5CUmfxmiXYLVJTqpoRjgfbeFAmdIuESV4LWj9
F532x24jMvky2kVv89iO3Arils09Ol7KvmP/dlPWbHJPXN6GlRuyMePK/N5M22R1oKEWXBWd3mrQ
MOFTh0lL4vLl3AT40sK0ZQuYb4+F3laDoG5n7IeIaWkXgBqTC5pMo8plf9c0AM0+yF9H4puhLy0j
BwgiHpdd72ovUuTDl2aBgzgBHGbqSBKvi6FM/gbq5sSUw4jClk2Ms3eA5UR38rwYebmSn7KChJ3s
zJcuehfi3Q5dO/3IsEvJuquiPqCCbU51SE8rwWQUy+K+JSUKGpdt36dX0jhLy/J+sJKkqCCT3AAy
IZNg6Giz1fA7csx2K3cWVAU83iC2Oo/PPkLBSjbDAnfP3d0XMzw2kPpkc5hALYdUMRxhf4FJmkiW
fPVUO3JfWUxJmjDgrwhFC1z4mpKytvT6r2tRBxsjMXJE2UKJq8A30KmzTb64f+syxbuezHY9au6S
PH+p+OzTe4lg71UkQZtVY55NnXl5nlGphrDXFo1tJ4mbGofgefqjfC5xV+yUGDrROPWRauZ9Q3yK
+YQaIEuvuHxORTfVDsvYcmKRRhXSHskZfJSM8gxMn2SB4qnNhoT+G2pPT3y+5yIPGYFHos/0gAP4
esqklyHq3ujV+kglgPS7NC03o+7HkXrtC1vOgnZbHQJ93FG/QfT/3i7Mrm4iXeNrYD8zgvyxIoBd
PJAXCCLSjaaLD0FQa1AsswEC3btzVDuWkoAxEU0v9JftsOLhV/jJJ9DCsio9/i1Zaaow8FQa7dOa
gVD5sqRdldkgH+Zu1F3lTzUrtXHODT8OPJoinDxi0bg1OPaQYFWgHyqMID3bS68fyoVPEgZ35EOm
4Lr81sc1raOqOjBaBvC/iLv8yP+J9Dd6yl7RSXWe2Y3tPFR57dkXoWBsAh4VCGfb3vhH2yZ9StXU
dZxsdKAyqNcnWffxOFWdTTB99EjIyOxLHtjPm99bheSoA2y70sxbeLe4TLzcnchVXAkgRep8Z25o
G241wWMbg+AanbwkInLwvTYLq41IOlQ6zMIHg0m4X6ej+BOUwJxGQWZvuFCixtVQn/YFXReYwJQk
lppTItut/t7Y7pr+sWye0wWV62hez5SFadOeiiwTJmCcMtaNwb7MssoajbMz+30Zi8nAmdPB14dO
1Xa0a7LI/c15Bgo3tsj67PLvO/xBCwto2Z4rM3jeO4WmvOzBFnLOD0lKiIhKRb5MOP+2vCOPTlrf
t/xtiZkcxIPwARbqnm/w1QI2oiAtlAjAjGBhJjlKZchTjblnPDbcX4t/m2bZioJFh/jMeBo6+HbL
DlgZQ/iJ9cjgAyJQK2LtOpI71Zq4m5iVIGB+Ri2HUll/o5jdefU1R5VEfg6Si1ReKrG7fiIbEwDD
DxBBC0qCavrUbOGXdnto0ABZB9zWAf4hYQfZ0z5Eq6wSSfg5c1xsHNjw0jBYzMtZZJyCQuJLnU58
jlK9RTdPVr5g0KiITJnuPM5G1wUIDzb43NQmNRFYvDDmhHhZgclbj+gDU0+YXHmuVBkSkSxHriwI
Tfh0X52JTKUOdjRWx9hZjtlOldWx0mRKxSENpmsrumYQBIBNFoerZEL+ntYLD8xLEYgfztdbcAE/
0VnUz3s1rQRjzJ56ooa16uRM7HA6o/QRzgAA8X8YHdKJQq9xYx0+laVHfAqB3seW7E8cnuNwDMax
o2Mg4y+JZ910v42hZwVohLM8JGJPM9pWKKLWyTCkgcOdro2c6WWVbueR3lJ20P6mKiBY+/AX4QAb
/CEKT3me+CWfqzFD6J3G3GtpC/Np/h3MmotZwf24hD2smGGWWOVTlvaYSc5utxXkpr23N02Ohrmm
ylPXMiXB+6dUMPFDDqbwvHIxVgsDrn1XjksDP9o3g12yyCHNzHQ3b1+5nGFKJ0T2qsk73gVcE7dg
5jwaG2K3UPq8hqG8R2SMn53Yw3v0wq/Tl9r9Esasew3BLwe1lnGiGAwGzia5cCTz201dX0bAawuX
wXJd3y3V8Jb6Zn624r+SwIhiQ0dkV+nTTmSfLlCzn7KzihycM4TdFsz/0KToYg1hXSQ/kMtOnkgO
sXdDm7TxHG9uGZfqbYoGE8/JM/MznceP6Y1s6f6d14NFl63542Azmn6DhqIsr9AGTlX9r959LQB8
a3kbwKZ0johaJS6G7s1qT89O/RSe2hJCz/xQmYaL4Lwl3GIGx/C3/E7/8N30d/i/2OxsZ13/rAsJ
0tV2a8fEUzbwCWIMbMkmLft6XvV5o+sEz3xvQk/ghfgLbs8TZZVjdgWcqAQ/z2MH3BOG+g5QHvgD
1hsu+JYN1VXwbY/sKkclUF0RlLl/oHKbAlCaRNtpohluNOj9j/ZaCkQAgiSjVyrUp8bJnVtD63uf
6W+2ezwUgL2hWajsr2kethNXUKe4Uf6LUHLP2rtb0Q9HEeg4+T0WUNd1VusVEj4wECJEBvyGnUY3
cvZQuUli6c4M/k/cBT8HoJBZxo3u/kOD9bAn+PtNkMb+sZUpmVEC84h64z7vly2YrpNesGBFzKAV
Lgtjqnx5mT2Zuvo9HRrKjDK4P2WBlZRmhawvOU0RsxdhK/u4aNW7fn7oTOpp+ut4O62w2a1WiFwD
vsWPorJrjqg8uSkKkhwkXyM9KBuawUMVe3r+0GFEOtwjDiOist5od3P/WeVCfExarkTDeHfTDSgf
K1bbLJBcQUgSU5jJBhtBAwmH8SoOP/qvdHbe6S9AkN1D4pWUuSU2+hYf83/jvXVRwxwCBZX4WJ1V
SEiSuycJ3aBapMjfLxwGNcIF6mNpW80PVkhN9apWgc+R+lv9i4ga6JaBr9wzLaf9N/FpPtu0gRuE
bjS21qpG2xcIh9Yorsb3uWr0zqRgI53cVSswwvw3VtP6Kx5DOsPypcx1X85cd2WkvsHVSdMVyuPd
PTSaWl4P1O+XrO5F6Kd4aaFaE1CAu7ONUievPtu/zzF3o9oeWg2MvahM3huAb9XyaJjq9jelsPbu
ootJuktp+uLwQVFSmwKvQ1lQuzjRZraf5difTwmimTtW0+fIK4Odus2UPPMdr7DjZ84af4igkdc/
GnhLmp3H/AWUUOhMxaZpKdNP/eBR8vxr526/IPFG98YXvdUqEJfso54q2Kdnno68f52j46RUwMD/
V3BajMUSzKZxYNucUSKb7/k4UotvvZhukzAGU/dt7LOCh0I/WGfSXc5fnypS3WbasetoNokox/+X
8sgue0JMXzcQEWjPzsSE8RfG6Eh5ZThaUJZupHvWq1F8eh3U6WcJFpLX/VyKYvfLaqihjF6LEDEV
rYSwlMmLsEbQiPj08taQBgj86/A7gQOMI/4Pk12uYmFS2VLgJl6NzMUgt+dhwr0FvADe6kl7Wgp5
2ciF7nsd5L5Ciy7OPLVd1yF/NGu+bN3pqFKiTSCEGLtAqs8kYLyVDYYXUT3lIydQPUAZmSd9YnLE
WTmBiiSHtPnkrW37rBS02hm2ayQHX/MgaHF0DRFRxA6+e0VtwxqGlJ0NFoqYYJBBMV0Am3uV/1aK
paPCwaCiqG6x8nnIAQ/ht5T/AHOTaKzy0bIDMkUteXhWpKyv3ACr9ZlDhOLUONjrRcZX+Ubwu5nx
34Lo3lb2wSKL7jwBHUDD/Psmh2tUrhczmsMK8tSzu01mqsoKQ45qZDlNTj3aD9IpLsWSGxc2+gVA
6PV/MvAP0NTTZfEd6J6HqmS049S/KOw4MsvcC+ACiSArnpJRuigj8EHe/9BAl/SUxAUkqL9H8zj9
YD74dSBTC5ZgQwiwjDnv6zLYB4MmY1G3KNH70AxVyxoJWzFjTAYjouKMwsCs5Uu73DN4IBh8/BZ9
7fhLINoRXYuDqMDmkWZR+1qN843BvVR5Cidt/i/GM5p8kQjyS4EK5kMClFfi7cAZefwXLk8nSxrC
FjPtEhn638oKhSKYFjECqmKaneI+SkCNOGlLrlIw2SO4AOJOBb4kgRnq5S2dK8KXr2rHZqP21rCl
/DV8DWhEA59iHdIUngRGGfXtC1w1Ql8bvHWHgScGGqyehl1TnPBj9JFZTZgLACYCqHoM45oAps5R
fz3ib63VmLEiFhwWOWMYC9Ce8u5qzy7/QHn3Tjh835mYxJiy9+EhOxHQSIteFU7axMUDyBv9LOTN
oOxjra47aUZk1C8sHbqqaalgcVMVZ6tmkPNAaXSAiMNTWUU4aQIM4wE66pvd7kJc5BKNiqjyBcBP
m/Tc2hcTkCbbdGDghb+BMA6LsWv3rFYE7T1z341+Nmve95Otp0HwEDrNfNb/B/fjG8LN/fsgsH8U
oQp75UE6C7kct9wI6oj2C0f1FsHtY0NkASi4UQCJzTtJbv4tbH/ENh/gcxUxztAiGLJb8NtoydJb
9bEeYCF3dMDdCDQlB79GCGvgoICIqOpSzQm58xT/3h2FBzunm4tNQaxerwY5SIa7SI6X8wdV2798
+dkVJTrztu1zgOvxsZ0P5mVKK6o6l1agynen//YGVcRqBa8TBmskd50Dl8WccyxO+rIlA4K8F47H
toQJNR9tYEdesRH6lSESYO/3Py2WjvQWqlYHTSgZNGqQoSPC0yeYcjZbuxjk1WHS6b9GFaujh8jV
6gAYNOURi1ikWdz0kxk79wC1AJn7YlD06mT0DLLvMdXUFlfFN0qs8f0QYFXIP//7sdDB5tFZJieT
Zhc8RCdHl0Zo0NRuS8WVSfUqPPruzNgRNKpy/jS8OZjmERCIt7u3xabCom9BK62muFwzuKpNwkq6
CtBR+y3RUZi0F7N5y6caMDiJW9eXD+mcDq48rFSwpXZ3kE8k077OfAWOx705gljER4z1oTS9uHg6
o3igdCmli2+JAXPvqpQk79hV5sXZFsxCrX2nr6xo/IlAQpLOmQeTg1YPLX8+w+jvbT/WQMRQNtri
NoPVZ6QHQ15hE7ThsOSI//zrSCXAkIKd4lci21eDHKV0zpWpRxNyv+gV8Sgl5dGcvPQOjGg+YfVQ
j87UeoPgwRaNHOcQgdWsxT/1BNBKLTW86duuvnWWi/dEq9gnpUdFCSPfDHCukC/P0wE1XhBo9CdS
UdqNg9xGpYkVXcJm38bAtER+EOKoJ6deFyQEAao51xpi/cl+iKcuD7TGvh9dL8osq5OLjNQkXCLX
qyAVPmJ2nzy0I4lm0lGkbpWhyd3/dsCq/qQP898DgaiidMD2T4QkWj8zy4YR+bFSlEAIA5VJcmiR
JbQ0USDXGNj7TQXKN5Reev7z2V8jo3xEiFtgbDMLQv6+QF5nK/3IJVQGqWK2JCiHKQ6G+2yMuDxI
CJfB2B1rHe/5DeLi9ZfX9aAx0sDrBXA8S7fuD9EW2cHOKhbfECvvmC6ekXdSBaM86Mf9bYMHabB3
DFWCoc5igh3kMxHKSkhdw9sJzaPSyDf36T1ZC5TtvOhftrHZBXipUVV+rC/ATVHEyCB7h0SlRyuj
7Ut56tFEt97IQGEHZTA+CdUK1qY1vp91UiZcneKobvytl8Y4cUJlQtGmG9JgizbBCM8inD1QNX0z
4Gto3pSJaVIU8dJWYbw5ycJgZRkwmgCeTmr2qxvptPsXqpIfkgOayfJ6J9FwPn5lSPCD2S0uI8k8
nXKMpFqeut4Xafgjj3TeGTFMNaNV0QFTzU9Lopq4L5H9Ha58oIdH4sjvNgXhZS+df5n+HwBP7WTF
J1iIX6SHnKOx5Oqegt1Wcy+FsGojbLch+dwaXUFm3toRoyIeiSDX4TsLII8wHuNjyC5NnRgte6Ry
sVEUY+RSFoiNHE1XLudS1VqZRn4lTSJtLiRKIn0HRmJWH9VHrIJVpSe6ggnd4d731PVJbyqkOaPY
Dy8iDNGhgtbIT5QMXP7iuQXKKe597N1mRzYgANMxOmn1xPmK9Wcih87Uu39ktnlz4LGIfgWua86c
YLlAYDKr4YaNUxSNPJIXROBkcqN5U1mg1Z1fluzjbHaYiaPpAVPPuL37jqrT2QBqJmuPWdjQyxMh
a2P/8/U8elCMCgvUCCj8SHIK9rGuURxYpdHW3A9rF6d1iLi/AQaog5I6sI8kdShGleMamw8i0CZn
0QFoOFHgVMAfpBmAxXA+kPXPZpT5qEzgY5ZzhHD9GdfB0v9FHjdPlnJEKoafjXgrhIAm2vURjotI
YExEn1kziP3/6GCcnfKpH9Q52Y+R4pbMK3T/S2RS/leb/hYZssxkzxGSn8hEyBsmxrfIckOz5vlA
aM11YXGhnRFfd1AHEtvsrKpBZWAIBT1NG7XgawS9j0Jxbo/wt6ttja+yEFaAINoNaigNLodNFRMH
H+F6EJArWOXZ+hobJ1KKMHs2ulGX9IuRenBkrM9QXZkqmGdqM8cP91wi5h8S0gxRdXt4qSVClbPL
puYkvufxDch+dWfym4FcUQOmGbnnP2KdO+oxQe+v24cgBGQv4BI/Osfy1YBg0OKmjHnUfefv214j
doR1uANfcLXsazPgQcfXVF3YzU0Afw1rm5cDkBsmnviLNkHIzQvNz9ljcDR/Atl2BlPXNP+FT4PH
VQ3/g6yXTHlnLasRIZUmAQb8jkWP/nqqMZ0NVCyuuBBxpRFGbKGLXYEyshejM68NyigG27KWOaUO
uiiUCZ9Q5K2mQGJY1GT2oljul4KOXnjCpR3rP1YQJ3BIqv7bHthwYofwaGf1UqmjdvqF63MvmQeA
GJvcvjwtMeGpm9DSLvA0/gq47xbSGEWcyXXAYu3OTAZdEB/V6qQduspaEBlM8Jpn8D7ELOzVMBhn
xB56xjqdGhNPojIVRvH8i15/9OEY4cits34BO5iJlCPLlNmIG1UT5mrwVyxTlt58b+5Q5nCGT+UI
u2Va4oumg0VyX8ppVawSLkPsoQFIV1Ty5ZbKe7Vr3p6Q5AW3sgALyZRgOmksAqxd42pBtvcG3e9v
3d7fdxZwlQ7mWvZI9XO5GH4eN3Vc26v86PxNEw2lLo6gRuojzgFDqGZ5LKyqZv1sJCyc9JgwNW7S
6yk3y2tqobOj4r/lThmJwPhLFH88LSBcWypoM1+OGP1YiKGEIyOW1YZdeFMIvDbYHv8tCwSPmx8d
3iEFy4jphpMlyeGmbIYyin3xvZDSI58FkZcjQ3vDr1ltp5XqsGLFHq8lSkTXCAAdb5yY0p7vKTTl
0sBPcw+wUEGXJyRkZG2kMl2IZ7PP8d3ZT33Kv+YR5wlhkWaVw0nvOTnvoF39ZL4tIqOkb5g2yxa3
PVQLgiB9uJXqnpwtoEXkBidvRJHAhbQwX7QgwcmwpZQTFnJsiLR6JV1z3Ag2h+hLCjX1s9liALdX
KT0zQy/N0ppE/q45Pq/VWpQLLRF1NRwHMg5AtAMvGUUQQ/ovKdI5RHPtmf72MVzZjiSjMPcdtF+V
5jKxSm/jxzdpw0KCefMj+TayUNSOe/jy58wLzUKpFy2jfFeNwbKiqoQXaQ9yf3GzFV1P3cQ0toB4
sZuJMPktdobangvBg82CXcjcKjl/ouzsGgmwZuJE3Sh+N942Vhj2BOEhSXdCm0i30HXPiva4uF43
dv564H0uLYipY4qhEBy/yfsfIarLD7QmdJ3wMEXoIr9i1Qcu7ouqYP8mirQOY8AtOyY3rxdI+tWi
oEbyevzrFa5NASytYbKkXfhJHNcu1e0BkrTVZxw5jF/j3eqCekb0yibvfcCpmBExSqH98wyJvVl7
QT6GXW8EAUAXJ212vtn1vy6bQNAnIdfaKD8CavTg2Vy1yLccxy6iLEb9H2yqo4lwbiFXkkI+NbzZ
3Q7wjixgKDZH4N14EYe6Z8XdsjgEM9bU+0j/GlV0gvw75+pqiY+9JK3p6De/quch7xXtNDk5Kloy
1rwaEjaGfDcU9rK0DTqgqaZW2SYYOv2FyHsKLX6d1OyJQVcd7f0STrw0obo8USV4QyA1G7FaHjqd
11R8Jm/5X4LWnh0jDip/eOPvIfH9f7r9+nuBMpZVyQNFYpOq9rhU69KnoU4jW4Kr+fQi64GrYvOw
YFm1XnzHyxpYP6TrpqhPV9RKTWvfnp5GqbPdRpgr96+IeZBINrFzD5FrV62EERt3TBw1TmuphUT7
O0QvWTuAIfS4c8lxUMvanstoEvNvi/klijiBy7ppIAgNTA7STLV0fAjLe7VkQsug8ze7if1zI9n7
Tft4S2nL64sliUznwIix4vYr8K3rcHBiVy5K5blHeLicwiITlo4EzKtuxdkFD/p7UpsCfjQpEtU1
T/1FaVZqU1TjWk7MwywH5bPs2TsXbNK8/PdEd/LwkO65ZdpEI+fFsP29kRYBmoWdDrHRNncw4pxn
CgvMHbROEwPmGGOIsMxx2fKjJ+KtJGZ6WQxNVUzsKYwRpDk3s/ObZCUsTQ2MYHOKn0GRuTYKawAD
iMVuWPAU8k0+p5Bgw0BjO09/fhaylKvF9Wz2EXswCs0nVB+1uZwmwVQ8zO4vTAp8bW3WKB9qm4za
8E2/Xu0+/e8B++2Ja5j0Cck+gs61ygCRKklKI0pv1Ma0+Hsf2RKy5ftO3Wadf3RPs3zqYdbMc81S
4+HAIYSBUhbEvne4WjZPZyxtw7/lk0uoQIr0E/WwzdjpKuc3xtf9JDSvCYBmr2wpyYPGIwQltyTQ
KYuIa0jtukRaVt/b+XFlTLQ3Z9Z36pu18+q8um5P8qX6mO9I7wR2JXekH0x0JH9rgj4eVLGjI8/i
SXPhfQLOMghQDxIZSR7MoXutWX4JAqEvTS5j+IudC/vk8yg6X1ii+dkQciyDj7Rqr92dmBpKWgKf
G1FG7gunF0H5TbCQUA71P6s6EqfmWGhRM9f+GlyxawyWet30W506qAAfvr6aOB86MxoFQ49BSHtJ
8Jk9wj5bHVsOe/G7u4D1RdENvVsn1XR0ZEMjlmPqA+Vd5gXDZxtq5yYwD87xOYBiM50Q54OyuzUK
zVcN3SJO3rxCoEJf8Fbmy4f7gg9MUVUS/qk44K/78eFfIL/1CkIOzORwGxJiU6qZV+mmCj7BPvjy
gVWZiMsHUd/1wrsDUy/ea/BkZaQtmS5JMHe4+o3j0WKuAXWvbAwlu5EygBqDwad9zwJp/aBdY5rY
fYTCGAO8j4ihbHew5/S+f7KOjvUijebdkFSSaYFV1jsafl5me6onMpC9HIkghhV7tnZreTHWtGMC
MN5/p1QTPEnH4BG69LwxssJmIZMxH1zGUUyo+10NwCDYhsMn5aFBk3nIgtBGMVSCQscDGTuMfVkO
g5BRIxhHKrOmq0sgx5oZtgD/TenJN/6TibKrMzGD6nG1n48+QoZSeXcnENItPdrZ8UlDAW1e5Mg7
n7Xmd/4V28YUa/6rfm8vxBLKRQ12Ag+rUWnRCAyBdgT6U/zNgAjWea5jyvECxwfY1GDsJ5Bu9CId
LS8y9K4zlpBTBX9p+BnIDAIPue4Zz+1SgktADqiYsut4D09hALTqcAutA9Ph4B8M1SXuupPzxF08
5gNkcDefPcb1Z3HvYgum0bxtB6jm6ytKUGg85barQisXwEJLCDIn0u0F7eBY9yNirBucR9CkOgd0
fSXxjLO7Thny+yoi6Y1ouexNYgx/pf2r900A2Lsw+u4CpgoNYf9YtcDAgIjxUCPPm8Ec2ya/5qF0
JF4zDaPAVYNGPMEhalhCvDzdXp8FoEb9L8gNtE5DCj0s//zVBurMAH+Cyfs/im0urTZWad5fsxZN
RcleT3/OTHpscq1eOqVKGl0TrSJh2IsYgDZbzhDG5qNZWUvjF7LyWexCUuGKk/Lmfd+bVvOsjyk3
+yWsKNIHmW54imW0ylLooxe87OX3PLyTrNf2d8zX5Yv/ialaO01f/lgoz04jzhgc7wC1NHjBBTSq
UOmAFFepy7iy3VHsIeUo3NKtPR1T1ialRo3cE7OPLpEBOXi39D8NfUtV0PgAaoKhhfPMVMRToJDR
zxOOoSh78feFVzRWCKg/0+vF3uJuY5B1tyzxcLC0sEvinm2RaXV0Eb/rSW6sG5e9hhTVYnXvcQcd
iL0m+G7Ux5Os1Bd9Zpjhs8/iEsFqE0aChLjiEYeWg3oYkYjAo0Kfn/QkkT2au67Nvc2tuOdlCdb8
XE03JmmxN+Ua6YVZflRiCZkllRokMspRsWJz7R4Z3JiTr78BYhivL93GWjP7sMOV+kk1sZ5RtxnN
7dpRuOTubwg+3IVE9wY70N7ejrqAVrlVPeJ64PFqWTQTTOzpm+uFHkLSvndyDho9Ij2ILpX2faO8
pDc2LFX60fKC4P07Bek33T+4ZvjUy1KAw5ZE0s/SyVMgIYIwBcIk/iCTQIcXHSrl3ZLY/Xc8GaQb
LmLsZhD/EmptJ36A2fmB7un6JNP5o+CviXmrMy/oadRhXfoFv0LNL0tbj/qnaRrJh+QOXS3mDD21
03j5kYXUsGpZecBARMF7h45mqqYMKtxIeSzzoy4TVqe73ohqhvYi6vN9vl99lOrjOl7AFOH9BsDR
XNzfwiGmdgCs1vSf0gHHpSZyVHK0HYF+mu3WCKqb8Ec/Iu+bNNGwraUYPlM608/MqCkKMHJ3xpdv
OCc1vJMBNU6sr6B3UkIMiPH09Ern/OuOpfW32y1IGOpwqYUWj3Hnnid9GiTDxdtR68PUeh/S1Err
kooki8Rrvk63PI7l7L67Xt4SP6zDyMeA6nK9MoB+ilROaK8VkGzSHXonJPET9yRPXZPaA+jMHt9d
1Rr/H3NUwHXIcffRpWfR76k2a7HVj3BveUZO9OD3jQCUpdkd1argu8cs8e8LPE8EGk3dvhpqq07e
nUddXucOMJkPspJa6g5Cj5OsxOCDl89fHJTVhakz3f1znIMJLcskX6Wfjr2RobtN2L1yeRTxGcZ5
mW1yJgQi4NxnwIvZoTvOlf8cfZyUW7GzzijTFKPilxcCkIp2vdGdHrYB61Se0em0PrERJ4d+tjrk
VOLbTcJWndr5cKH9fze9JM3vFhdItmoELzwHg3CdtZpNaD5XdUVWC0/X8AdGm6U/8Z2UPpZKIlBz
hML7oTDcrIUdz0rE/q4Lu+PXRIf2C0Ehvbxcnx00GAXx+ph8qFtA/mki4ws5sXFDfa0Y2FBO8ELO
JSsCxCpapLnIMeMA8es66ZQhGu8ELKuaeclnzOG32wl0zcr4jLbyhZ3qn4ehiziIh2FW4EB8YQFH
Wzq6bshjieLG6Dnk9RdRPNSxcaQ7Z6ADpYut3v+PSrRVpYr1olMGG0HCxshaVxdIwkStP6w6TkCc
N1xvppTBzqemSZwXOsHJ2UYYNrIZt3ob66wQ9zR82qazSWrVD9HIXEumH2i3RhdBWpMj1PpwC83i
xMMO1/QzS0l4/emnUiQgw/RkLK3UKqW0VEqyC1tWYnQFrNXAHrjTDxdCCvIzcpkiGM1ORo1ZPYel
1Q0XG3Jn1kn6qFW1aSq2ZbgrfUVC5XyRXZMZzAPZIXuoICaZClMOYwleO00wzh812wsJyFYSW87x
V/tE5WLQQ2qfp0Hcubi9rUrYP8jhLBhWnPTdgeInHAv2YSEA483Nk/PRMPv95WUN51DLQIvF7mAl
1gRpUw/hctj+QvWeS06lTpwEwQUP7q7UANXQOtZbX72VdIhR1H6nbvxP0Jxak6PJswLTMIzLGKcp
heFI2cIQRdDNpWQ60VusX/JePLfwf+6aFoQ5bTobF/EJi30NANVbmkCkgfrBrxVJkBGNc+y1KR3z
YIM58cnskEauBXk8YobdkhMbLBm+UBz2jbU8aTsvDlkCEt2UllVl/yGC7BdL/G0/mvH4xL1SzpIL
e5bhfcdM2JRrsaSrBmJLeV9eDLk8H8CDa1KWE/+1rGvc8vLRywgfRL1psE7dGoD28cDB8hKE9I/n
2avbH4nbrufGO1pS3D0iksrIdZO3whvLAMIw3nf9xB7bc674jPacmZb0Eb+Va2XyFYNRPzm+klin
MlwUBVWKCitOrF+LP7tGfeqFMF1H/nQcxI8rufa9ENs4NNqwXHqIiOjG14fVXdYAwJrKZuiw819u
iM7zhgOBs02nVl36L/IF9NQu5xiz4WYf3T1Pu0+rwiXP5mEUUBWiZA4jOqaRdI2stwelGq05LWrz
ViWzDYVikyhqw3faif0SbtgD4eUAUcICgVIouLbpCvCk4brVGB/20fQHOyBJNdY027WJjB2tza+r
OQFAuWnP08ssa2ThZ2YgUv3Q4jDCAiR15qvdegf/jQuz6hdv9zCCgZaElPOCXuiurrcjMK8IA3MB
4jghuO8zCUbQuQh8oildRiMcOHisLZa3VvQe2iubNKJBe4lUAq9Naf6S1ubZvYDn2xkJuXqOrkeC
SbtWSswiqrnk5RhKJsp48uTPMB3YPY/e1x/WQ2tRQU+ijPGf/q+b2B/adhEGacnbi64TLzkSLyZn
HgIhhL/KwEEiA41BPXokeiocDUus7SCfoGu04YMx1aAzHpSeZniwy46mPoxU8RcO2gnvnKeEssU7
xzBSMgDEWQb664/dHhEeW4BJPHftbDovpRr7rUWg4LEnIhnSnhVc9rNMjCpxbP3SKjQr46c1vI81
y5glZ/QhwVkyYXZ3aR9l4fADAcjyCrI3NJTED+lmyn6zGaABFRaOzOAfHxIta0MWDoHgk7LO524h
akLuJw/t0ZDwqKnfp7cciBZ9/SsPPRimc8hRjNpVigF1QimcGnJVd2ePNPVMvQFWBisL3BUak22s
a6GcnjbEuDO1sLoqZWxXXR3Px6sDZ2q426v9lLwSbux386jz10EvVgEZO/KHRWxEeVSYZ5bZK2id
eAyf4I/DO+QIO7/NoSxwlrZk0QngK7+uykV8000qHMDiIGjoCIpB4/7+oQwXDkw8heia6tK/gZDi
ytd3EL89may6BVsiqY+m8e9HM/msxpN07PI7vnXZOI3VoyvQT3ButDzhpFQ1ODZHced89i3Itqs4
NjryU8r90hJKJIUMZZvdL558cDfjlx8CJVsysDaH30K3OvLZ7kB3TAf3JcMt2qZ+BNrINh0tdTPh
O1oHnvUGmZDNSm4467qkAgkpzHXWrhlyfCMeD5/f8ANsfqpukvAwhYXjHkxyNW/FTqzRgowtngBm
KPByJ5HM8KdxneTdoUJIkBWD1ZUUXm3OcbR13vciHfbUfyT0JGYutDul22T+C+fLcD3dPVHqeBDc
YpaeI6+/rKFDTZIGmRz1+smQQX5/8+rWDS4IJkTw5k2ijIkzvYg0yl5dTE3soBw13WoU3bWksVDb
XbDZriLkT3rRmkyRCp05zpQMXggXhTqG8x2SyFOrn75ic/HZGc0LXWNufpw0VPijvHfncx+BQX9H
xoCvvervORBbOpfuNFr7WwMqqdwJvL4xgWz3e8hS+VBofMLaRN60K8vsomYIjYINSHIjZgImsUft
sWPEEjqQFkuOlBzvW1kDeZm2/fH7lVZggMd8b005VYdf3Cp4YuGnNQJCXzrho2Um5ncVSjFCADMM
9jKNVDHUCVwmkckgzsFRKDUtyrNzWDh/a+ekk/QRy45sdfGUSG1n+t87Nrb8kPvrS78XbiCdoQ6E
dXDibr6/tWG4QBlM3L0Pv/EPm63NoXb6ZrK+tQHR8+AwB1s+LyPRc6vk/UFYjVzrVP7FItL9E66A
z0yepT1NN7v50SX8RNVPiVBYwEQKRyQQxRqPoHqxLu/enctwZYH92oxQ2t0VxaNfFLEQFKIUliPi
5xunL2nu7AkCJZc7MC4JNW6o30aTt9dri9sRK8xABhY2vSI840enT0wdTtmGaGpsJhPoLkBtC1Wl
UnzRPJirPCbZen/O1rSKkBXCZvMqH/sr3bU9tnWWcrLUutSD8GsQkgUR817kJ333sxerhToK7HkK
ddaQ25+junRahkstGvk7xbFHXzRlhnPopGy0r388vV2dkZWecIB9eEb6x62h1U0udmkemvpswRVV
Tio+lNzvGUDycQqVQ//FT+OElz+DWI/2biE5j5+w6LfCMav9vR4lLKHq91GGTrrzUC+x44Q89xql
COM8fpdREEskupMRLUmjHlZg0F8fOX9o4s4t23rtDb4tKuNuai8ECV/S21NrJoAQyEsyOiBihkvS
r5RJNiMuEAGGqVzr4oeER3JbUAGoDsjVgOzBvE6AKsagwONr4YxNY9kmn89BpdQD13k/cof9Te0Z
DygpDCNsM9oNbK+/42nlfJ7NqZ/2Tcp6lPRGfsUerrY81iL5CQefkEmKnkvCSnN702eh+H6w407o
mU5Xk0dT6lR85Wc7Oe2OMKNbqPhpqgMWkgTjNLnZV6xQbQ0QsLCei9k83U6RLhX1M1v52eyEwJYF
v1xQ2XE21kqcjE7bikWm2DLvi3bdr06VLxhU9xL+fdu6UXy4pUY5zzy7rl29jTNWRiJGlzCsVbpV
y9IPppN2UJFJAN5au0m+q+GBkde2mxbcBn8EpTDZVFfdjBUTCaPFk4jNsHWFwOEz7c+1i1oLPnOB
k6O0JKWSOO5GdCBgwUYe9a2XSzkGWh0qc3JYpPQ3Kl4P8oExkszaUz0HEVnNHhOtn9yD+kptp7Np
bpi8+V1bmITMWx5safN7o8ymbaILw05mmP6uJQpcoph4UQDN9Fg4YUsdEnEe3IlaE/xuZbrU/FOh
duC4aVhAqXU6Zw0W6SxgLJu/o4NCiJYa6vM8DHNFN/6SavPzTFNwZ91A3/MFgMR/n/ztUt3OKrTZ
5cuaI1KfPusqD8Nd3dDaLYYmvsEnWr1rjL9/JGCysXJmLivymtKMklYfkiT0mjIUpbZuuZ3HIPzL
To5KBmZktiy21FiTUXrfbLaxfCHYAvRwtGyaLELhuw0NCVvuQi84RcUTx38h7kitBvWzQajk7AK1
4tLyOadwSwOq3LJMLxvsBe7nqku1QfkqtZJfkRWPzFRQtIVoSzAcg2jfmbpO7GByBNHCjO7h2fza
eYvYBiveD8potHZd3LSDHwEbZTKqgLFaVFaaXNaeSZrJCkNUzFZdvDSK4AI+S9M4SEk/488YkWGg
r1W0FwT0qCphzFsGDvroz88TDYer/LuuFplkVBbFOdRGv2wuLc+jXN/zVIJ0wubQjObYeixvkG0u
ZVy5LZHh1fpMuY4lV0P+8gyxAH047dOhq+Sr3GUK5gjfQJSX/Bk7il8cRpyAcctZgRCCzzs5bM+z
L8UD75g8qlPSBaFgjXDdrj4C4UgC9ULDxNnYr4DqHBhqHFOvnBeI8z4gUwjS5gZvD+H4ymQkg+A8
Mcimzulx//bLHC1YI4DB5uApf04eDLMeF3f6KUh8Qygo44gYTB816L9a3qxSWMleI91w1BpjQQPF
2NsmD9FIC2UArsaopmJAHv+cgbrBCmp6MeuWhU76hHgCcYdKdI5411I+p6Ujq1ZRAramGBwW7RjL
DcY+DLmH9yTzIz47JtexE8F5ZbiYmTNxk+U2FjJHo9P4XdmlBfqBO0mF1oN4UYTCIYVI9+gW5Qkm
Uu51JhlGEsBmROxLSNEmZ3/5mnqCtRsROhUaWpP+p5rgakcfETJ3aCkogjxM9i8IeUjBqXKQ5NZz
Ghse9H2eOAs5ggy4o9jJTztoqxEBdKwyw9J5tPSqVgBqkNj2O1UqsRDs7UCkPrWJ1Jo6GHDj2iuW
cEEarOTRDg0KNJoKWJF1wvCcc/9qqRU3srANFgVBmvK4ftWe1pn0/xB8iwAPHUCA4TW5GI7Q5DBm
LG2kAghhFEhkbI1IStiPKGKGpMiiGUk7Asm5086c2NMWDuSKxRQFBfSbNDyy/wzEOIjNXuNYCAvP
q+HFTBbcbXwfJJaaO/yqFYNiYzT+xFwQsfe4Mq0dvuJkw4e7ugbxYqvviQ4yC95xLxvy3AgViFOy
rqXGczLg38yugvgwP5KwU7cIb0KH8ar8NrhuCAx6gm9e+ckDoqbVMV9zcGKNFsM9RE53s/DCtAFn
rYcuvjBxVc8TMhduut2OQ2i4Aia+D2wptNfAx6KaB8D1y41YbtIxDn9aEee3jW7zH2micl+Xkdkk
24kHlS2Xxrc+VN3Oy9/POszttQ2A1BZTRCnUGtce1mHv90lhxRsLA6IO5EfkKem2b67OHZibvDRv
HjUnZ/0QsVCZjP+XC6P5rLr+ceMMiVXQuDQURSzrXDlY7KX79mC5qqprAcc7B3YEYdpZvVR9DSl1
AnDOh5wY3Aw0JaZZiWqh3JC8Ovbm6pkcTK7qjT0U8Vdp5vVv4udmjLvZGp5glyMPCu3arNeoh0Wg
S6pczHWkfO7aNyk8QS2nCRtTmgTGGFWmluRu4sl6s+cb/9bil4L91mM9pSpiU4fKnOhvDfmBpeG4
HY04LbAkdLM8QGZc/bpqXHS2SNwnucKyl1WmqHobFihQ5IahAvo/vATfcBrrqSjnX1kNGt2RvXVN
UaVN0dDhDMOCwkAHv1dpRmIq5DpH0NasdIyqdSALZURZb8Wiq0cSmdbRgZwHOxqh+HWXxSz9k31m
XrmESahxO+y0bfNiu2QDUC+ranDGd3tWR6qZkVteO9Q+6t7FDoX6+M7+ZWVvSvzkTJTZDPrF6BS8
1WBtB0iaoe7melbwKZZ95xxFzHOi+2DqAXb5ZVZggSQ1R/wmRL0V8FuVDT39DZlbTufhDoS66BBu
QxXKNWUzaqqkXQ8pVJ2MMVuacDEjnrkwZDjFsXVxntw0JgDkXd5zaajajU89L1E6b/gtAYlokEiY
dH65aNrfAFWwig+5qj8fSzmPGptoD4GBQY66QzZm+33FnNpiUyi6JxEBbxuJySpOLxB+HsPlcvyC
LJKwWkxOD++kMdDF5mS8DLIheiVmEgYgmitmssyAwwePckx1e9yvOfoSS0tNH6WSRZLPyx9NGoX6
wSoT7co40HXnLxPJguQb30cRF7+1id+U1iFi5IF6d21OdCAGy2sUUqsYI7qNtuDUm7x7CgwLN6ih
rSnab12z8aQySvQakX6Z361kCO/IZrsJwXoWOn8GeBTktcqM6LfVta0UjCMglhYHvohYVFBYtY4d
03hYJKRMRMwKOEfpD+NYeAYwsNvDI+FzY3KT77Gmt328+zg1xqI9pC9iucJYNlYAHtym/F8uxixc
ym37/O9i2PaFrsMrk34M8H0mVIJN4+2HGmHwxMWcsfYXIElSuACUIbLgdasJrd2b04RmuKfyGJJg
Ise7YeQIl+XVTT+qfY2RfqWNpJJajsSJRD+7iPWrUUtcCf0ulbPJsV38ZBxBsgv/Slzn9dd6xjnM
Skt94ktp57VNPluQqpZeZWPCUjrOiKb67wesy6YjueZvbxoeKxiVFlC2hYjkVDZ9ybybELzYfqz+
gLIsYvweQ9Qi5jk9fezTWO3xW+b8W/0j1dpwiYamRp4FlyKux406BcGK3AqJA7ZdLuyhShQRgiDI
mZyafeXe+9NieucmCW1XkXYMdxyWaFw6NCXKWFtXrMNUZHXDADpCRzJZ8mE+7TJz0HhLwGbJGGnR
mp6qMvrPaGZ533UTiO6TkyadEzqbHpZtQ316s8kjCA8+L3jqGjMalF49W59n1DyMkQYdiPQIFHD/
3FYYi/1QjfaQHYDXDptYvU8QpvvzbI5HFHPfJCkMW9DeETwipUF8bnjmS2t7B1JYp1YKxcJG0krl
6ISjNYYpxyaQ+cqmEvPXaW4MrW0ja4U10GqGrct+McBJUOUq21CrxkQERldLUbDC6HqtPFPanPi8
SHYuh7vq3INPumgQ1g6E6+zDp2jnFJdPMDSLAiiU3ffbjNG8wdekR13sriEC7UitoahgAWWitpPr
THZJEm+1UHEUmzTSkwg5DXZ+Hffqdu1/TG06V5M9+G2ES27TyERgYpt8EmJqlyWxp/Gg5Ui+8+cH
uT4wJLQdwRaKb8yD0RbWRSjGlWZnLZbXRmyUrWOrp9/akes/HXqlqI66tj09GZg6zU4UYU/ZPCv6
QzpX/sWDO3hIhtYUNhjsCfHoNbH7a1VNg6wmyUDL/NMXAVu7u0bF66CDqVjiLxxu8qzbynoNBt/8
QT2fnhzkyFUwBHZa0Dbd2nHEa9Ny8cOSynlcCE06+11mCAKF9znbZvHvSB+MOK5+AyghzCyZNbKu
O3Fb5WbS/HoqNedoEDwt2DsMo+6ZY9dseCjByXA853kSe0yvLpp6xVyqccSrqdhZ1qJVxmrenkFZ
HLPW+7rjh9TRtrMDkrIg5vvyqe+LQK1NTD54oHBVDQcUAI86b6S4MAkZq47JKpsUQPqyYDxPAK94
sOUGemPXYF0xjosNGPTkUuswVu0sDNC0yva1dnOPKuZHI+JSP5Wnntl1TPM1MQB8ELV9MIZ/cumJ
K5Z7oKlc3uI8Z6BtERnOrkGICl/US9RyblCFkUCtoDdQNFKBNmqfUqEq/274GltjX0OiGU2b5aMV
qAhLNiHXmgo39cMg/rkRZG+DjQNE5ClyWoB65xMPmNylvO93mpa+VdPS6jMGMqjl+68WQwYrnsto
0Lf2IPHBkwAbzvRSOrEhspI0Nwz8F9CAy3rJjWKFJvNP4L9M7QFGy31cCJ8HNBOi70JHxK3MmuRb
7B/rhzEROGSFcufJbrdcUKfL3H/hX+S8D31svt4Po/oZe4byD0stqML4inCk9Wi/B7qTnmniMtHC
dJHbgMumTSpKZMf5X1BmeqGF+ZfAvuHA8GXuhd91TfjdPy/zxcri6DhqQdORC77ruOHKRZDqqNT5
Wn3+saNVmBAV5WTFOVF0gpJGejmGU8fBQT8wV3RFoRcrjs3RLaY0qaK4c9f+8UHQQEiNk3m6bbZ9
naviiP0rGntP5kRBse+NpkU68HPg3zeric3bfWOv+ngQWUySQ4VXiB1dcffDwm7kO4lh+m1OkDc+
GWfkrHJlUp2BcUXReXemToQJLRpdPPsLLVzWdTSvMzmTXNkGCIpomsMYHTPrGf5CuPIlWjNnoOs4
BnzbHg+t4N/XJZ/CH+w39LGDu7Ds7mo/4tp8dg8RcT30wFgot88gCifoZZJVPxPXNKFo6JdUDXYG
3CL/rcMJ5DUulHlqWxn3m6ZMU+r28CHDxyKzAHnfYDa0zpf1TSoMDZMSM3FsPbfWEtIWIxDCQwwp
zFkitMtBE8Asz9Pf7Ipk4AY1lEobFTXsvZgehh7/LJ4V7YhHz1XE7ycxVcRMIephfSrUrNRXS5+G
pP+JCCcYSOMlnlB3kFJHW6o5XwplxX1xwVdxiG6KIjHF3jUYJ1+5cdoCmFhdXSg/eaxCcYTYgqVD
i83xGHeRQf7jxkTr1iIEwsUuFauikgkh5SB+RWGOa3E6hYEH7MtiSpP7b2n3Z+5N5bEgZiibUTcc
WW/58I5ezLy44FBxMd+8WADk60r3I+J0f5qyAyhrNoVcb2WYHJAUJ4atgsfQYbCU8ZR/GqMsI7kZ
JUvn/UY99em6Mcquegyc8yMldhv4RKlcCrPwORFQ153Y2LlSgcI6dUk9BJx12HYaVdA6zf4DujA3
T8YxO6Cuu7s880+0FztC30WYUT4vRggc1KO4y7NIgsKV3qE/xa3WB0EdVmwwQ64NXMTLl63ORS+A
sdQUG2gnve8zxKV1ociKIcdiMX/20KYhPqzXrVLIcpUWo2RjT+uz+pXcPfN7lUJpuvQwgyllixoA
Z9YOYlXbgEq0VjCpWf0MHgHu8+ku90AmUKYfWCoHnrzlXisbMhlD6LNhu+VNDaMgi6blikh/KDGW
O4YILN6xFA6L63msVCSfDsuglJPl1Ab/uyIzbmPz+JJj+DA8XLkn/+8Yzb58fH4Ur+qKCd8jGXaU
doUn5CE+tjEECR/hEk2jzVEd8El4I0pMBW3HyNE/Vm68uUlfHOimqxBIwZ41eoZfRHd1WfShOGs5
ZNlLmSaNGxRb69dZqACj45xjRD2ZCNkQDfEApPhjA9IIpeNqwUz/VNvoVtPRFyn7yBxmbHcJ91M0
ANm1CSCFHkXSKEw6KqMe/Ny1uCVGqS1theOWyPxlKE1nmPTJG2+elqYzy1uckAJlKDd2w2YBZCal
/4FL420PKaSzoD/qMYtX/hhJwYSYBIe7pa3jCXes3/HOOXjP9vN/0SzGbnKSo5JzIIHFsaMCDh3U
AhjWK0uGHZiaucBHHFLyrgl9DLaqcraBnimp4SUwR/e7Y5Gr84XGbLloYWEpYICpFDsa8HeP2l6H
VbuZM3MjVhW9F2ed9VefXcPwG8fBLaGpuC2BZCO6WEsC8C/m9ALEPWcrn3Gw6mRst28+3yBlJYzv
lDgluAmpsIeK64PX4TaeNn8mrs8K3JMmdYQj0XSxNgdq1Wh8h81d+hlua5bi0Qm+Css0n8UBPqCA
UPYsJAEQ2m4BLd8C7Mk1VNvoUDXsdCQzKo6GwAPN4LbjRnXBwri0gIwh+Y4rlrFxjhXTXpHJ1Anx
B9ootW5Z77f7/8aczekH/g2tujo0iBGSMymeOoCvVfx/mY02VplvHvHGGvDz2plGACTc0jMWHDxT
/CHfBU3HBVbef6WsxSu7dPRncg78UCbyOLirNqdxN3BvTElX9dq0fK0VCfPu7cjnpzaeleMWRDcb
O1P6Y5fyU8zSkYvJ1tT6ocW3j8n+BCD0SNwe10CMdb1uuKeHXlLaoukd3jGIxPlS7tZB4/W5n83y
bUvAHLPhQpxYWdXiLvFOJmBkSNcHNYdNcdPidc9YLh/TeuUWWDH8EyHARWobnV9nH9GqhsHOSsdg
EGhL46xhypCDOf3AHKiMASsb3FokRfRqdKVTrzd3mekc5Kd7GNN/bKUJWojl+eNjh4G+WNNlu23e
tAsk6wKo8wbBCiSWfuiJTgzDxIcWDoF7Aqe7/uMDGBFMmB19ly4MtzfgCUfNEeTQYSnBh6SsCyfb
0J6BUMu2fmhbLINZF+TN5GynoTqu4kKSFROHdIxF0xRejGWP00Us8fN0PSvtquYwS3wMev1z//nC
E7rboEz0DCEFMR3t+r6q7It0l1hynPpnycvnVxutjRddzJGUDfa8zfsGhn6UBQjGKjHfShexA0rg
zcrH2+W/zRALibIULlV932PlwO1p+zTDYLYp7NjTm383wvLzfwpnA8XeCeswVq8p110Vm5qLI83h
TzSM5G02YmcIWiGS86HuH+aMxU8p7Ahhms3cWxJGmn0jrfJi7DDySAbpGJ94KvX8zyXWKbBAF82R
jorFWK+PyfHzBIqvRqN0UgC+cjNkqKUh+82fsPjNSgTO4Qvm9xyFp6IZu5XJUUROiNbq/IZPDgC1
rAAkbdQLCSmxMocbtlGRCMygTd2ZV6rSZTdzPDLJu/Wj1befVqYKBYnNAJGyGLviJqOymhbFRgPE
bQII+hWFQPKzzVjNRsd5R2sEosgpYzg7ej32wLqvj7QWrMoa6PagKkm3FZfr7Lt4eQK9WhW0/ZUn
3GNYVqMuTsijzeh8xs3t9URAY0l/QxVii2i0Tax8qk1Y5f6tpPtKJeqtl5mOI9Fx+PZVur/wnUqX
PzCyD7eWlsXe6cUmbrt5MQqsooAShKTpyxpaAC8RV4YBN3weyOOpzNqA++FEuwvf9qoo26axeCSX
HjOrrqBHMExmSoZXvg6gJ7TzeBLl+7oD+2xMGiKihQiqWqiYaxo4O3ctv7XSubBW2aJAsskTE2vd
aJJSORslivpqr3yth4qyXC6KIc3pitNEbA/r8vcQW1lCxriGwS2OLQuq4PDYijkQQtco8pgGN8r9
Xx4WVuDJ/SKSWQS4Gp1P2E8nVtBhsNEH5AsiQjkggTSTkTmX/AUQSZ97xgv4kK1nJtRjq71OYMQJ
s1gyh2DfzJdokXKAWThC8PJk2YjyBRq4u5lwg5Bzb9at3EomAw2TR2IkTC9JiGFlPOTIfK5m4SZV
WKiqvuHEr1dt1GK9HTFXcyeiCAM3++5JfhaBwqwMPTw41y2Uc+D5Jn0AWnCclem+YRsrNh+Nwplm
LJ82zINNTC4MxpLVCYtWctdOhexgvH7+QsLTFc0WzzkVfXmsSiPDAf5ZN/z+Xk043L03RUwlJ6bI
BJfNIVnRY9uZjODfhwTBl8AMFsuh8CU4T/+edUpui5fsKXrx+p10z8MvoLSzOdAjMgbB37kQ1agN
7FFuq4nseNuuAZIi4OH3KqQJehfJSc8NBl/5MziCgDmof3Aq2KpgaCMyQeOLQrORfTqMA5B6MOnB
Wzn9ilVhqnI6CbYTYH8ywoT3jOkBi/GQ7rUJgibdeP+iEqNXeEW49CtNn7TzTwaGasAUySIKL+eL
2ms81nHNaeCugxUUQZ86XrGnq3CPtLdSwm18GggK9K29nhaod6e+X+Z+pTvZ8UBzvBJz4l1PjS9b
X1p2SCqhu7GeLX2peqxlVGtdas3W0O022BYi2ppUVq1OFhxqQiM/ECXtqmUH1m+26o/kVTkO4Tlj
eipHud+Jt/pH1w7KJ7yRsanjIjzb5uk1akqRepUKavP21R//7jesIwF9Zz+o4KuhUuNzhe8R9tGt
7En0+oQyDsdmZluL6LMG4zykOLCaRIoem2ZmLOZri4USBUjwNnELcOqZ13BPfC5n+PwOwZauaXAT
e849Jyc1ZgBHGB50awJ6ERdh54xitZj//9YkvXdYidkBPr/jp4PbHNHnC/V9I2Ml73Uw/qXJ6h0o
aiF0PhxDfS0wU6elGX12iSTKnaP4/dEtojrF0TaGZPSAnRlcP9FRGREW/CoGEYRkjtHyx8luKrPa
X+mf+jXzTipI7VSbZg34pyjehOL+JvHgdSzppXsJ7dMN8MdJCLoIC9zMQC/k3kK5SdGYLr63ZLPr
DppJjvLZAwcnpkVP+HkyVCMsZFkgT8t2IxyNZMBC3iZwoA31w996S55WMegJkfTlLtRiEBah0rwC
aVTIfkQC+l3xwXLhhZsWbkBow6IibqsxnR1pI7WK/o7tfEwQDJGko+g9J90wKE9llyVdsVxi/R2c
Kk0MMeUbl7MN1GDyUXNlIWFxSfLY39rG4yuZ8+Jx++h/kmFwubtMFmy5dGmX2Jabx2MDD6gKkeqY
f/K76CfXcORJ8X5GnQyJ0CFRMU3gx1cnpeVtgJxYsbzG6XBNhcdYvv8J2fWYHthaInANPj7bnGyr
EEHqzKJBMep/VpOWq5XUPMtOiq2JgrerEiOjXc54+mNbqXBmWM07KWL6SnpOWoh5Py8OzoFZXAj6
JeT0/JsXffjRyEloVBisJDIHvLh5tXdWh6GDAfkR2aeHUDyvjAEIaMTZHzikTqeUDHguluriYKf4
6znVqeCkxvQJdYFZK0uAHep+SoDLgBb8BGyEyAaMvbB9n6xfVR91LiHc76NpZ/7MKAFw47LD5Ev3
1YlC5WjcTqxeCTIxtECAxq+40NdoXeRwL1DO7kyu46qGslwIMklqS+kgx0B/7QKCfCQlD0x9xlCR
IeU/huVq+xcDmbF7kfXlba5Ty1eDDa0CQRd46mUhaT68f3Ud/KFAADnwt+TXXYviB6v9Nnlll4Z3
Q1i6toyb6nTP3zyNKEHjxoJ2STV0S3p0wtFOEok6i29rIBG7gMfXFQkQZ+wAdjWWdxvg5viBxRtK
vkvdtCAW2m8l4w15jEX872aBoMtg7k26IxFq3sUKMs/BI/XOJolRZUsxHcqKW2nZOqow7gnN/gT9
SLYnOvQtxRpZfKfHU4qgghnCqfOOYk6ZZC9m4qxUn1D2Zyb5iKap1wo4iBanNJ/xVTNS0Se4iFLh
eMTjNei09QTNcPfcXqS8sy1i1TrpyUZ3ZPyauZgFpDfjQBVS9w22aG55MCid+ciGZ42P1NcpfJrS
mTLE3CKfiLGZh/LnBPmaRVpY0YUNY5Rsb+YKQlhjY5Zv2LrFTM/8edJFqcGNGV9HTSO3YGEQ8OD1
iQyRO+9cgvzfL82dz749j2bTrLLOsEhrk+0wQ230oZ3CG8YmbOYLI8xzwQfVzL/JuU+X8bdvl92r
4wKUQwlshKgGkFYKD8gvzWi1hnOjcoZd15BFbh/MmgyEZiuZMcZUQfQDpAHntAC2h9th5C7mRbp7
JhPYWCpWFTBwgeD/8w/fmnLBF20VABQZVXfgCeikGQKP40Bb3RQtYsqhdJ77Vu/zPODLIRg5b0rL
koabr6/X/DT1QcoO9uY69vf9urB+y0uLxzVyZ5FyZnNlmktkjNYnfOqHc0wxPJJTknKAdYUhPWgX
hLI7fYz83OGiysgkraqJkvQQYP9Q6xkLwdE8nz/9eYoXXzY151e4Y/u0Sg5ZLTTjS5UeWcG/5wuQ
geIltQe+KFeyEMQ+yH0IWeNYzY2SO18yZgdNRh8+pSGWtLgkT+71iJjHjdtCiYv7VJf3vF7GPCn6
TbJbMKZRLHVi59SYDjMd4DhiO9IvbnI2LsXiyKCsETnmX53aTy+mSoKWo4BRVSkszQ18YsJgiu7n
zUAKVDychCY3+51RKhM99QHbauyqAnwdG9M7Jy0fUp/9mbB8U32rj+vb7oGxx7Fbegpsg/Ee/gfM
ZP4MxjsbMg3EztgLy07HLuQxB+tSH1fX1z7IcWQBn4ISKOHbdW1jZze7sD+i8B+8WSFponah9A/q
xi8v78PxGhncjDz3FwSo11A9iRtonEztTu7YcAH8DBffzzbaISmlvnjprmcFB8ZZqbAJvd0oeHBr
19C20P7HSFPiXLrwbI8XCdY/++ikDeM3i8lm7y4TekM841hqKGbfa/I4dsqbVqcFAvfTiBrJTWIP
m4VWyCAPKOt1uozs+VpFy5boIUJx3zwPGEl6Z5Bu/WY/I/ccmhY3z4W81Oud/O7z39+RjnnY77U3
Ytd7jq+8Jp/EcKaKzibTZQATfNyk8Qan1wY5g3Q+bgfS9MPLx0YVPk7UrSbCvHyc5KBx6JxKhmeu
FirTB0BNO36pDey/47wOarj9CdLj1sF8k7NO2DcUY6mUxf0p/kpwZ/h/UNB65aIbF/B951nGtXlm
ELvQm2kEmk9QHgERfkjwBr3+atXN1wMecuoxY6ECrAS2X83PUJi1XvENvJKTZQWa1SA/K6nHIjPQ
0wcIoUiRaxBgTLPgvI5GIoCPH2Pqk/vmPJr7s/HG80d6tLFMaHCxHmWydupvQ8I1CCqt4EzhY2xN
32Al+MxuMV7ReVBDDuBvPmgrnQk0lKHm+W3C+KslDTI/2rAkHuYFdSVUBVcs0FZr/L/dThs3NGsY
lbbSDmBp3hTeBdCxMvTsOzOdODQuEjjlTOfjTTNa3QQ11t663ac43KKsKRd2PCZQNSo1maYks3rc
8s6HZbiFDQJyjYRZHzlGSGXT2ScSJrZEyXa/Jw9AjlCLdQNeQpK/Z4tBcQfD6enfRf/AJL3VOql8
ow6v/kdjEGKXiqec35RlpNLJJWag4yaM6EQDVpfzzMApHfbZ/G48zczEvJz4erBDq96Wa/6haKb+
suZwoI5/9p20FanInq0eyNhEUUZxZ7usNzctgc8tvtOqMZkU22LRHYMhPDmoYBwmE84GPyzsYgZl
HeoWBFeChqrNFs4Ak+/AawpxYd5qSnEzN6a2t3F/ebis/DjuFQaT98SgkDeG56tNSCdziESOfSvQ
i6yEe9036g6i8iVdchFrWJlZC1WH9sxx/ucPFv432LkAuuH+eCQHpo53Sd1CeK0fGLGFiSbnRy5P
adXRGfoqNXL6GeOQsYkh4DsKz7bFd+fs6G8x52CertUR4CsFu5C/IigdDEcnFmbzHmJRHiMCi+zw
xoY0UP1Zat8uS+t+PQQiK91rdCgPFu+D+C6Y3CTeaNP6gJTQymX+r2f1GHLyZUNU653MPFlRqKCY
uzYuRrr/gCHyLs86QO0T+Xq0kcvgZa4nifk/HDiL1N3Ij2iKhpd96R2Ec7/EoKzb/V6JPozJw/OQ
UHAsTyNxFFlNbZ5AyToBF/mBbeIyhg2bM0ICqBL6SOR/Xb9OoXU3qe2nPgwKPHU55iFstuicCFPa
7EpuTzyCGyPwc1ULO45CvBusM10w2KePL6Q2jVVnKQHQzUIncWqjMfeIINqPhJRXQV8rSuUqxeAz
SNVgVQ8LegFxgSuHUr2SJn8GMgL8zEc5nXIdJoTkHFzBDRVs6q/4+0TBsu1UCKH+aNrSffFxyQ7/
xGM7xlwYZO4i6q8BJYgpCYdgf5IdRwGf0bUyCLhk+hHfWc8C/cR6zU6o6ma7rlqiTYejDbXmI6FY
wMwze1CTgncYPAezBti6ISy2JiiC8nqOwF5DZrOYVsGyMm5abZydYzm1xI1Nhp62fx1VXrfh5u89
5hTKhGXJxum1D/oFNmVIjxIBaRmjoVIXUOua/xU8USKqajx3YD5rRwQvjA327TyZucGXO8wAildy
/1MVuQdM5lkzIrZS7Oelch0uiz9CRIvB/jhOfpBQ3TXwlZLUetEQACtMhE8WL9yweR81cWZQ8bF1
qQo6X70KgJKv9ecVHQDvGOlFGyX5ubbEGlmwqgcK0rgMa5gZfG2LBKYqSEB0TrQe75D53Meux0uA
ri5idm/N0Njp+PFG6IxKhijL1vh0vQcYydXbB54nSLk7yEmHtDeNAs3b//pLp3ODXq/AuJzdxGA+
0C1UPROczZgg7xaU+WsWkQOzde/VJF58ED+TLgQOwIMigmqcEThfKh1Agrd6Wp/IGJHGtQHr9UzC
DK2jDLiQh6iRGwkncyLAxaYTqjAvceDdYTb+Mhz4IReMSktpHnqEMJAWhWMyjQTuKuMRjzUwMnY4
qHYj0NiDzGnFEpXhDoZX/80JPd1LJn+FxU6rilq6cAHXrQqn3Qwi5W7UL8SRtk9ft9gQMNeKoFZv
IbUYsDpMsTinmE/xcFxuBcMlbhjF+xk1UN3SpOBQFcGxcuuClSJRmmk8XQmgSLh01zxAzA0AqxPA
8VUxWf1WSv/vSgXjN2+JydlIAzxRNmi2dEMS1+LBvcoyiRlmuzE2CkgKqiD4xaR7s7vN4ZLCh/74
tCDj8Mn2odQ81TWxCVFmzXxnGoPwkuWC/zcLZlhBWAf4qqC601XWqiSa5Ns3okAQ3kpibU80xnss
2F9vyUognQUUY3bRusZSWbBP06p6tMkB6lveqnbqxtIzVGQrMFC/0QS2DOd8nySPWKMamFITjhwg
saAg0s0vb6TfoUKhoriAHPJjJbmxMFz6gbO6c3xzHyyqEXnCjHG0pXo3tp8dhvfSa2loZyrlNd0G
ChduuQ5Yw38wBbGn7uZdzzaZrihzxzJQj8RucTwE8McIkCHR9Kg3HPE0lLRUTFdQ4YkY9dnVnok3
OInJcYpGm+XVXRCHxGMs5AhvAamhs4HFYI8syIpiee1o6pFR/dBmgGFLkf1rGGlQGZYAwjcn+Uz0
NGLMcnv0pWPldeNWS99MExFBJbZ5JF8GR5jsFlorouK4E61imdyoknHbWJnkpi52zlqMqvlb+G1T
qemCy4mgur8/HgMSZDX8lT8m7bXCAyAAsm41N78b8eYW9/j8sC1wzGwqB07ILGrxrv0HAilhVrZb
EMyp+o3K+hvWCsbzpWr7Dk/rBX+MtboVzwUiy9lHupVnm3h3XqA1jt9YxWf3rCmlhClOiNFj+Cdo
D2sWzwKy2lcYy2WcWFGSN5QpMaurwyb+1XD0hdxagcE2uWmUwCJPwUb/d9vlJjdX1zg6esUTJHsL
UVZM6PugjW13F/Y57Ai6T8jfZBp5lYfx4GsP1gouzxkMLZfXLcH5k3OFoxKPSD3zSgRyjmfYXOnY
/tK/XQo/AFx195GKJIOA0e8c0oPJBfe4ow6ropjk4gHlE80zKIjr7W+NRtRfp1nF8O0Wj7+W8LKb
xChK/hev9lJavvEYCxDFMs+/Z3hf7340vFFezsxeiTMhhPTrlLh8JPN4TwJ648QvDQtgzU6+bFT2
WAFOwQKECUFAd5lIcXk7Yuo1yjlYMx4uFWxHG2jmMf6F4RwgXtM3VbTg7vc4OWtcDe3ngpgdXSxT
sOGBTp/7os4Jb1gOP8M57o4Yf0MGCuR6xJnxNyA8GZ3saquYpJgrPrn/K9+ge38ZhFO5x7cC9PWj
qgvSEm4nw/fRmzP48M/62x28kGpnudIjuleSjKa5t83PIEvKVlEXXs+0XWJPZe7PjDiHYiFw+0iD
EF0/9bn1HTjQcZQf7r9GBgm9cQ4+fwansNTdFp2jr+QUMSOjczi0u71e5LAXccrGcSn8gzrzzIJm
h7XOOFfnRDOTm/xIs+ZXqhIWViQOjQpLukFDXjJ2b5G0yRJ0NJmMyoytO2zmSuGae257Ek+0Sg4b
dd734kgb7S89P8DFcDUBLUdzCl6J0e2SavGhThKBk9c+ozRpBGcuGNWQ3FY0ssb1k9SwVnFBXXYL
BkWHd+ebK7lzXPfgL/7ZgJPjqaYKLS5Ae8UJ2Vpbd6/31k5oQX0mBnhJMrx3xKg/62/mCQLkfNnf
Xqsk2+bFteXUT7LqEJQjH6aIkcVoR9XxST6xE53WrBCsQsDAbAy2yvinOBLv0QggZsvdFTuFi5eC
caHuEJPURPy60nOqAP28Rh4lc0NXgOQLcD8XM3QHe80ETvwEJYL1BhkyRrHBbIIVkHvTNRHAdT8P
Omk/zKPh8Orbx/z/K4CAEN7AJ8c/o31M/uG51hk+Xn0VC9GpT+rAgYAhjOoK2B174mNiCjmp1LxG
qfvKrT/HvQNUE5PR4uBiyuz3nzIF9KAL/cj+8VUjTOMCS+lkyKLQvOljOs26C7dU6zpIPjqcB7ni
4BK7z+0AQQcOs82xMqLAl3z5jg2HXnGojQTTuePLJeqtF4O2KKScw7iHMQeSkfMPih4OAq15Wd4E
uo3tXpng4XmAt5DNIwKy+NqSd3RPbuiu7wNdFbJV9gDOVipvz+nLmCZYDJRQIufMZDyjxN2spkJ2
Rs99CorR9NKOqhJJeuWCwBzOMHxVU25nL2hLMEwjatqGm3vuGbcl/p5BdSmqIjZ+s3AyLVmWxKjw
Ao1TJTa9mLf8F4hX0c3kyQdnUib8mVWXiR3uKw68mOEKjjrW7fSOk8li3pbfB2K1w9nSjkMvwBmN
isHw+Qau5ZQfeosBxde74Rae60ZSGqI8WCm7Ee0iP71cahEJCsMwS0yToo+8LXH2HtDAK9HTFgUF
8ozWysmEcrCJndA4JG77WxNqM0R9Pi+/rqu4rqUiMg9PDTcEdyVswWwcOnwgdkwGeDUjgf/jly1o
RP+PUpAbQHo8elHjp/V6mi8h2CiyWN6vRI3mak2K/ptRJqIkZ5Ln94HFnnZYkA5NTwTxYITZbCTM
QWRi2bYdpPHqVlHyF4zw4HJitPXcfsm4L6ifFjcFoSsvYCBCklQGSria4bn5qxK+tS1a7/tsAXvN
aRkOm345fySpEEAqNT6NIoi27Ol0T+YE1QoK6gJDBVudQsdb/OZb7oumiX4lTTOJBBNd7ROVj4Cb
jjHMa4zQok7kE/nP8vPdtBAc+rp5vaATeVXOI/gAF7N9vhHDKse/OTfsUZ8q+u5JnKabMFP/WsuP
2GMZKMv5PiVqBZvzMO9NewBpl7+JmDgNyqHcvTPXCuWRNHEvtPTSwo6Oo5v0mSsGTT+m+RpkFKxf
WMleAhvBWwmzBtjMZwJ+96Mk+I/olIuiNSJHxvbG7wTywmUGVocYK5nZJKiV0OgT2fvMz1qUFrEG
+VZNPvp/1WtURc6DWDuTPl46Rp2l58bcG85EnoteO64RXKi5TH3SvOE6X3w2ghmL0/3O+uZ6OxYA
bxES67pitOCBV2vkRrEteub1gefv6jMf1ORFugKQ3XY4T3YNERBmdiHn6H71lkoGKsjuUuqGg7IB
h9pe6h7368tlFPFtvs+NexUyiXRy5V3pGx1pTNvY//SbJfMvxLgMD/8rH2gYETyYocKgL3S+8LeI
gYqSD+yLduByS+SKNh+/vx7nLqnWINsuLEy8G4Xm7/UxwMfJfPcMK5O+9pFo3MB1kKcLeEqG0T0z
Wau8nfLpKpYJQ4EHJMgDY6xdPJytJ/fJZI2cg3JvMK9V++ilb6Te47EdJkyH04PrZjYeN/MpanhQ
6/kIjJ5O9wt8xQhZqh3YEA6019evCCqn5IGgYds5FAinZ89EB13Rwe9qHJyTMQMhi9CMkaEOdGF2
bxAN7OK1wNknYpooVFiJLKRcDzuL2NNhOrQ1/Gc6Q9IDuEOBRP1t4JY4T1FbndbcZ3ywWoukpaUh
e0gQ82cgZ9MrCiPNa5slKCI0Fh/rWMQ0TyaFVvaDHiAWCE/L3uFfx9UCDWR0JCRP7zgA6XiAKo3L
x1uGWVxY1ecJJSrnj28u5uDWzugllBn/twOcBrTaJk2mrJ3V+N6W+woNtRJPciOY2rAZYQ3SbL+P
2vMqsSm0ZBdNUM5xOC3cb/oRuVR2bhyO72b1acKnUzRu4PxbMygkffJ4Q8/XZZOfdaiOl20cOY71
0ANXylCToQJe5INI5P1yi1E4acYKsMt3agzyp4dT2oZvAjmKdJDYtNvZYaHYYRDrMeeGCN1dRjkH
F2WKtYaQNZHpYzTu1Vsou40P1uKQA05XX77va6yx6glg6pFwXqd4mBWFujLb8zlg5/ZvgDH3oW0X
wr0s6kypOXojmXixs/GO6AIEukeebouFh07tZOADyu3IWvJEtMln+ff8blotvqTsp28eeYr/nWQV
qovitY2AgOIlEKFCI7UmZeVKIxCyLYkJ4Gb8kBIw8JrMYIK+paHuYyLU7DQlsY/+VNisolHd/MqA
hKA7NmfO3VJiybCj7eyrc1o6M6qUBSO9+QEqBnoASjBxYk4Xkw607HDGFIhgL5ulds4tnzzJatg/
9SA/JDLeNEbzq4YDP+nnSz0GQMSqkPxgqfUJQdIXvPePz/uKQCs1mr4P3792bukLs0k5/YzjeDY4
4mN7YxkBO5RdIeERsyNG8Ocs1R1lBzESv92Z2jcDekra9zVv39msnQpmV50RmbG2YsEjirvKPPnQ
K8EI7etByVzQgic92wSa7m6X/N7LGQWDNgrZIMVjIKDYF7DikP1b2EKK0lnxL/qll57mKJ1LvJXB
OJ6J/MWM7zWpUQTwKV9gCDiQiviRX3TQXOWQLrfpaPSuRP9Io/iJg9nNAUHHLKmSLRGpMhF8xVg2
iTl1C/QMLVrqGDDYnimcyQyRt0x6ofPCN9M5a2Y2Nv91HXM9eVScizhkBUpm04TY6TI1o6oSkHGd
fwFu5MakzDwFDJE0P4jB9KGe20/tuEcq7yWUgeDv+XqN2/Gg75Q5J6uW3894zBOsA1Eilhs0Qqaj
0j1h0Zl+0s1brpgio94xXVkjy+ojtHdAm9/iigq3+w7y9XGx6FioYOTBuwMRmVozKhzQHGj40Qgw
7UeBBSQBeRo1pFuK/od4rBvDncRTAFbC5z+jseo03dTlG2Bx3bsQpX8I8AtSgDb+Kc2dPFkTj/DD
dW9n2LVFVu290L7fXXuJktAmA/qhvD+SJVudSYuWDGmu3HV/zxsH4J81UEBj++awEEWQsmTgsBDr
T65LVYOP+/AOvAbVPsUIvrlQd6ArjyK+qi9qOBZ69btGKprudGHvJgjL01IHCjr3kMPlxvlv6Vtp
CHqLmJWykWDCdMwS8SBWv4LpeIGl7U1g5BUJL50w9ui1WryWpBnnAW+3rVdIlqRtcrwT6dgVmvnh
5lkiykrtI2/XCJiKNqnZ4ODMGjeKOpkNMyiBCMQ++ad/47gh9JVDNGg+i3fuCw0E0ZJgmiHwYpIz
ogL5pPWlUS/24LLCUQlGx3pyP73WmwU0IR85ZA7atHCEbrfHRxLVoT7pxfWZftaxAqPigv7JMU81
mxX7ezTEC2f8WZhafv0H9PrIuiXSr015uZA61bXPxmwRJaWO728BiskSu9qL84pnhjAv2QPARY0I
/GyO/MdFOyudF7AUAE/VTZBjJrmGqtcNQxRTmqMcFP8wmmzyczYaZY/nhFQf2Y3dMOBX0x0no/ah
SAQ9x5BUR0YSejIj3V8JiMKHRQV8oE9s8yYBXM5R6W47jIl4xi13+/VJmNmtuDqnBIs1xKGOWg46
2Asn9n6+tCuVdSNZ6foaXfkn+I3OHrjaJJrF6k41f+zNDrz3AKVkzgxD4Pbax6h0/D8azSSjLUqY
km/3hIgBqaw6E3wAzJSZvro+z5ZBQAoMjFTKeWtnoRYcOO23vks9JnUlX8ppjeoUKSdHFWUDfO72
5aX9pfLE0m+JoyNk4/1eKCjT48k0GrJettwdU2whgYX3bVzPfV0v6i21a0B7SVRMdOYmbiNPk8Bu
OICuPapwazZErZn7vf/8vaLdD1o6UHDScQJSTnMCUgWdqjWmCCqHjMXFIpZa7dv8tuX64TGcGls9
urMYRFUITUaZPleYTmV0m16quuDjxobgAPSkIjkwtV0TTsDnbZhQa25vj5OPrD+QwrtIX125Cpbq
URjMgU20uDyNbEQud89XEStYqYkfQDPM8gRcL5Z6VZCVhsyzstDUnbVwKgVXyyjqmQMEOlWwS6Ql
xukRH1LSdkOXcW5pFZuDtLUUMor2XljSqGjKIdXF4JP9/UhRh05dr6xJwRuSrBrPQUY8GuL8I7Up
4GaSHnbDiT5QOCwtxsv7AbNNhkHQNsw0pl1GUHI20+jDM1c+WddYZAQtvEzr6LUqjQlld5BOo4S7
7h3QqWMJ8iq88+OP3vskMURHh92iEBoWUPTCb1P5WS086ptEAtS8gWOqF3GoiOP181k7yHjNb1vB
+B8JsABQsXSShVfs0JCWEAC5WURE9YyejtFHYytOPYOQiC+Rjfzn3jmLUJUATCLHkqYedM04Do/9
hYPHLTWf5X3KeOFei/InHV/FZHTuqaPmibbYNwWhupEKk9ep6FIaX0FccrV4cDzH5z+xkWPryoT8
OdtpmyAk0Dau8wVYULLWxRsa0Dm8POQ/A8sVzVMGSzkfq5JnXwD7nKH8UXthF+x9d5hzy0eAtTex
O2V+uqGl+nX0OwJwNy8TU8gwpn669gYR3ghbPmGcKr/liDWrYn5glIzdhsjvWjWpWkD/YJhzOJnv
XiTnKF3L2ZZ5hdUyI/LTDnxnOmT2seHlisKI0VNNSxOuAp7EOiLvjpFeeOwa4k84qrr57wiwmM+X
gJ8SginFRoajBYvMINjuhDNBBIzgUSw5dS7MA5SaosCFgXqb4BM7iCsORDcg2bYfj4gntOM+seZ+
pbmqXoClMiTutyBieTqQrrQS/sWi8xz1QlT4TWSvIM3VfvfbwolXu0NsHRV76mVr3IjoB9VIm06M
+xJ0j7ievWTwa6ZGEayJtxTmrfAbtLmF/NFjNtfz7tfPMJKmQnGK/BZSVDfWA7+CD2G5dGW4/vlu
v0jgWOQuqi21t4nbn7bdBAU+E9JGeVsBRUlLuvIzkd1r6QH3YPn/G2YnrI4YB0kdOkaasuZ3eL2n
KArjXrIillvUep48lIiteboMB3l40zATHefgQ48Ek3PljJHAeGI5oHmqqJ4F2n5whPHqBNcKZA5P
20sKQT0Qz78Qp2V8wTO3xcKchxsW6gZ2WBnr3SNv4231kO9OFW+aj37xPc4AwjBZHZpKvniyw2hW
gJAQ+Uer2D8kxNuW4Ea6KyK2YUa4tfOFONPkHJqhUpIuSvEpitGkOLOLVssp/IQz58O6Ki3p/A+v
um5eMNUo+gLp07wPxCOpI8kvqGngB+BfOnXt0DwcZ9g+3JlBa2HdHCIQ89KAcxbr++CeXT2eweEH
DgL20OpehHny+lNcBVS8Tz99duKRS7kvvem9JDcs0/B3hNh6rHkXZgAG4H7xemTwYqBva0QrqYKO
/JUy3dKVXtlFBxAbVIZmFfH/N7HWD7xL098dF1pLMrF4539rPmBzKgm4FlcskUOqra5yD/lzNAiO
3WZkJM3WZ1PfX2gkYyQGjNn9N31ZeE0RcUgt9mtPCyodA/VZZY6DWK/UX22V5K0y6cCUpnXGOZwA
sBpL2h2TWU/ptyXC00hp/1ONaYrA7qLPxqI9k90iuv123Mteoqi4diABc4p0AtmTBW5kmoRYg3CR
mtoRwc7xSaavsKJz2+8HSE3ESvjYJIsINRitqVd7utNiThM8WcO5Rc9wd92KIMQ8eHVPPFanAYL/
w2gzBA6FPBhdITEXxc3hkBLwg9PHXHxEDtrpDGds5sMk7ueh9uJazxBZHaHve0g0X09dOwZUxOCz
92sIhxbhH0dGsBRAxC/IMvkXkaSpQICAhp+zOG96yrn+0DPVWO39Oj4blMuu+SXT2Hi6In3rTEIe
M/9rJL2TSC9dlSDg1UwiTs9pZXDp9WZhYBkHYemSwOowKPYy2gpLN3AAHBbB89G1ddZhbZV4gd+9
MDBWMmXN0D22YiEHAHB7VwvW3EdChC6k1u6c6tUUnIesk5+SaZ/yWP3oszOTXWT8C5LoHUFPK1id
6fe94VgDqv8e0BB6MrulwdBkw7n886DD3XysGwskIIEkVkKSxBGlM0ckr1zlsdsPsoPpIqxpJv0l
0rpy5jgn1NqYkDb/axZUwT+s7gzSk6R0lu7731SMHBXt/XspAV2UTDlezTEHTYWrq+XoFxQEt4hs
UEfQzsA1Y0DesfaYysEXqrtu2G3637NTIXIfGckQ3NMMo56HqIXFSsiDhUSzIbEXVq9VmXcG9baP
K928jt9gSF2OtHX7LuWdlJgt1/dbonNxpJRMspnzSzzrNe7ptoN2ifJ8M0qh3RnwIs9xfm13jfdW
4yqM6mtcXZXSqA32p9i7uObWSzjAZ704D9j4wdQ5GKGMk58s/bR3Xsfpo+7Alhzzm6wzEZpzHfbO
XlIVp6RG1BXlEiGHsYKOt3ERkbd8pOzmDIntajpNLoKPXsTe9H1wYgcK2RwwfEHCHYXwaTmAAPcr
SyLSmFJQiM3FluK2H5KN0FU6cCMsXDHBNvycYGoarPT7h7UodX2QhM7R8sAe3jzIcdFjgX2M/uIs
c7DWePOP5VT06hYcVi3oUOQ4G4XwDOCCM3scuCIbTW1un65kHzk+aFYOj7vryjuTXwEnTvjONd0D
8OD3tqfdGCyJT+mzsKUUVaFm9LQ4Ta0XLM7q/HTj9H3A2SJ8UrJKOgAavJWBS8GMufMT3svWJZBx
kVqjzU5wOh5sNNdnuieNny/lQ2nAfcMfC2HzYFFozTQhLCXfPsOuf99fjOgs4NIAyCq62yGwnaM8
FbPVI0YDLjyq7LqtDrNAPLXT3PeItVU4xyQZc/w9jMRU87XWCRgLwl/HNzJHvp5ExPUIR/RvloQz
6xHqGynx1t7Kufw6Rjw65VgQCndap2dVrDj5Sj9mf00sN4p8Jxf8+i+mRgiePcC2gAbgkTjc9F9Q
ACQUtkVVB2C03mneeKsyDkWb49Fvq3VgDHl3up07yxaXkxN6wyvQUeZXuFKVA33O0JLvwsJNY9nF
lbNmKnAPNJaDDUamGVaYraEeMykn01tZh331Ra7umBnoOvzuYPPVAT4BK2luve8C90fhTMP3mAmc
kCku6u6CfgMp0hyvib+4dqvT3rkTTlPcHue+lka+z5Vlz57486EhrOxgmoj8LQt313W3k8uPPSLs
dmwtPINp3qll+9eev64UhUCsAb/gCDBFymLMDm04MotPuF11P1dbOmZTXT3BdzFzK5MvSJMuwrqL
vdMVU+RUi01OJHxW3hi5gwLjOTht9Vi3fLzOf6mgkbI9kifOHx5c0Qk+EE+zy6u1A9CLng9uFsw/
M2IN4bXAmfYk2jSMv6uQN9q1ZKf++XkluX1lzUNbQEGVYlmjYV0Sl6rU3Hy6cVNnZERwJMyFz0dk
2NJLXmyU+4oTJ/vWxZJPnML0w4jf1Ns7GqOjSU9RpmPGNy1tx+Gx6/eARhl8YcQdjt+0t8a/wZKv
Ez61jOvRoYBMjywq6dYWKw9GdwZyerdrRFhxnDT/O+08nD1EmBm+U8Tpv0PyG30aucGj1Ol6y4xV
NaO51UgnuvqMsgABgz0Lxy6kP8bsJrG3J+fulk7seyaYYzP3TIed2QaCLVFMdBIMM+MZzVbnzvgB
ojAx5Cr0s9c7rVcHijGucruELov7XjaHhXguolp6/XsmWG7h+yRCWYCHATR7+RGHkMsScrKd9iZO
8S6cGenTbxL8BXmnmJip/wxzV7J/KlTMDF1LS1SH5ldeS5affVVDgglNKnpsuftNmnNBQd0xRs6P
mhcMp4CcNc7KVAhBISGY6ODRIWjLkc8cZ8hWCMa0sg9jSpK8qooZXd+0yXoaUMQFq2DvQeohqrJE
kc387KZq4NjzPVkfMrDNhsmnwwYP22NesSVq2mya7+jwU1wGTnxFeiIfZN8e0aF59lXQDR28GCop
Sbg9oO5YVfNgNw/CaV4coaIr3yXpItK0kMhCUVcqvaiRaPaXIDmsQYQqMAVVi4twdHk7oyFYx4w/
vCe+mA76+U8CX7xbr8txad67E16m2IjJ+LaQ9TaZ3LF5ApX6dp35Wq4pHVfNiE3Bo2TjKdFD15gB
AGyMJwND+E+wefjLa3uqBPhqnWg4QEAG/gnWnREwY2ww1pv67L0rPWdTsoZ1Im6bfOWt/XT7WozW
rcIM5LRtc0s9bAfkftkV1Sbq4H/+FshPB7FbbbZqwrLAhp4rXzVXIElinuC0kJYD+yQYLVuCHQsy
tTZcf7KNgJ3mZbJfGs5Nh8Hwc4N719ZblmEdtr/RvFMeDiU+vMfkc+jMTisKbfm0nWp677+HY4/Y
/EiNSYfSGLw/zTGH6xcLiv5ZbAWOXVG7ObTbPkE1OUSIZFPOR+CcDrWkvgFgj3gVGK15mXrdeUiA
W1ar26UbHYSxqkFrXiB5GByP81h6dKf6Wzuo5XgXqYwgSU8S5DkTswaA9JoFq49ozXsNzaM+V0eQ
FnQaaf9XeinztHISEJKGp6MHJ88xc70KzG4ow/2wt6/9+PBf0V262bJ5jz9AYLDh5w1xgo9Xu7mE
cFd7WjsFkYjiZ/1oJl7KrTr1rmgylNKATDnp0z8oENxKaX4hHYh4d5C/WasIV0QitIP19Aw36eui
C98/6HDoPYfic1xAsZuwN2RHibBbMZxFlcmq8SA+tRSssa4Ip51mUYMqFVtBMj1NpwVOv7lX2Pms
xb3vAnlNeokFnztLN2XB/4sFTDQnzTR9/vVkAhfUEwUCMgYZ7poel+uYhyQ5iR2EHLd2LwNM0mB/
ZVdd+dai6VQLTleSc3cFlAZDn4t0B4xmNRk6volOaQ3VBSpDGfzQsO7Ev7bo/TiwUk2jA1/OMKbH
2kdPtT0cYmJaQCCGe6if097AckpO+n5jTXNq9LSSMK9L3RI0cPqEGXadQUSCJ5gLoBwruZTBRRLY
dzzBMeC8SOj6JEhdPbKBskeItb482zMsT87VztfwBG6i+LdmSdqivqCLuXhwotTJTZoIc8tlCkau
o1ZfyUc/d3uRzMe8mpoDDS7es5qZNuXRzf1o8rrcn7OXeHYJBWGJ/WT45W8XBwhpNX/YNp27mmft
5sLScnnzMrjNRq69H+jEATjGPaci7a1gq48ec/EtC4f9HwOQbWYjGBbkFGuK78oEH2lHhvz7YElG
lLuOPG6oX/0zwSUGa5+RbgHiUjzfxP9b7oV+kgmbtIxMB2OxVC9LsVttf5VibiktMVLcAl7tq3C9
Sicbs+akOFZ2lW/5XYu+xwmm9xcy4nsLm2VyTIMUWFCgJLx1HrYLGKNSH8uJtAn+sfqVrVTMVQQl
DSZ/FYu15J4mdXqIVqFWKznh81w+XzH8RyTVGc4zUmr/WbJ+kgx/PXD4Q+6mm04zkaT+GS7cUj2f
1cxZfuEh1D8zwIAVzq//eMwPCjiQhEBh94OLhByKh7qyrFzP25Kh/O6DIhpM6VooGKTOqDR+uU5+
UnWWzCnNKqnBU/SATzugoCURGV3gNLkq42twsSskLlnm75x963b4VS6P30BkMu3F0udJG69dUiNq
92nLpQswW5yYCc6NoIOkXqIm50VNLM73k2UF45YhHMXW6iuBOlsWRILcW1OoBxKyrwI+WMZ/r+yL
2VdSGzSL2mrmRCytuSotLpzX4w0jYe7SgTiOWTXDn879FcNA+IMTJT/iIeyxtwKuOWWDrer5DbF3
fuMIjgLnfbnQFPLOHjfssxIKza2oaEDrhdadlaSzQQYjp9eH/6DAtJdyTC4QL93ADM1TC/8YzWNO
Sjrb21kZxr7JhwZkvBrsEfDlD3V6WXidvBXx/w0qAxx+4eFpYYATJQqL7BvmdUxypFCvU1iDI58a
Fv3u7tZcei8FZN9WwdsgC1nHa0ZHn0pAaSTCYFL1a273s8eWpieT+3KaAFpJjCP81ERXuOph15kj
0XlV9N6ZuWmvq8GlNcWCsMcfMaWRdHFAddYd8QqYlDI6eT7dXNcFrv/LlWR9UvwPvKDuXmYBc54E
aYQsy7i0mf5bF83sENy+ceSkfY2IQdSVAJcr3AIIYEL8Qi952X8sFLSI0kyGmRnzkxdM4HazzTuO
EsHdXu5yoUk6uhJ8eZi4ecftye19xbDZimzf8MGRRGAvSAo0JdfM6QBNvR+MKNfRW249EopTkshA
wcePmFQspRXEalpM3WD6fow3GigPB1NXT44oUMt1ruea2Omiy9O1yj8T63CzV7/3HBO6oZyO2mM4
1c4fxJKJQKavkQABjo0ZcKFgT2htfWDnJF3ldKTFF3baDhZlTyRwqZNfYJ2BKau7HW0hjWqUs2xI
7HZ+lAL4X0MDYrpGVrDpQNgwP6qlpPuB0Njs2wUHuK+l/RZHBZw4du7zKwIRddYJCV4V/Dhm5Gox
7ZvhwFMIfYThRwvgKDyrhut+pLY0DyHgu0BVAjVpik1MjPtJ0POgWShVzX4FVH1X7k3aQGjPLt4F
f2rU+11NaYQgSfmBG2e2/2HNc93yIvkoEXYKzjxrs2pqJSIiA1gxa0xCk9e5F3xBSaRqcU4rd9+B
/Ea9m54Ei5XMmWXa1Jq54XlqrhOKgUWCzucgEnY75OFTyH6Wwr8CMcyIsHL6JtjaYyKTOfYsrM5Z
AOYUMWT3WFl/xdRN0uIQiT8fAWVMDWGGezPco/jC1X1i76fX6PLWh7JMnuF1i6DKPinyThNWI9oz
ip8iv1MRGWWcl/GhXXk71QgO4aBXmGDEgdTvm8vnbCqtaAfviKysepNqPztQwrKwvyvQdVUYcAuw
27arbF3eBAwTLnvWLY10kj/VGQCvuFNsFOMfGiZvP6IM7YYwW9MztBgwEKTxPnNwhFOPUkoYDX4L
PbMOcm38sHEAoqiZndNLIO2bt58VghUMmuKbYODWMWAwtvs+LCWtvcXjj0qLkHJ6LPZBCzV0Y9x9
f/JyscPFAOt8z2IuFQCLqh2d+1zGJS6TEUl6/EU0/iIW6Ai0sdYirtMNuihEv79UCL/mBZVk55Jo
xUhwyP54GTXjVod3XuAwp5/Byrd34hmXWyBiisbqU7RFjc/zCu97xd9e9pZnfXkatzcnfTd0lwrU
/Ck+Ih3f1l//9bXxfcWJ9n4GZzwi3wdv7iSBq+LQKm/21PqnncQUfg9WwjD5AlIW1R4w/3fXKUCD
m0R1llkAlZPUvYyK5IU5j5a9j8u6r7rn2a+rXjmlAD+q2gy2GnMUPzbTIikWRlIHinf/Zb6km+V6
jevZPIv/aTshqceI/ocjcjWbhniMJnFOeng81e/811reb1Yl8+2MT8HVVA75xGkLfilu1GMxjAOf
zRoEyUCxfgENkqr1Dr/HKzP+LtztqZ86G2yNcXg/mKG5R4tqE7Vxp8QXI/y+J+HJQBVSdE2dnTRY
IWr7oKCr/y5W4SNAGtjfl8A7HuqYyzUQGbIlPkSvreeAdQfYJ053HrQdZG5P5UMNjMjazuaZ9jzu
NJyOoA4KGaZCY80NH+wquzzS7QMYW9XgxD6PA6zAHu6Cqqp8upCpDzUn/Dw+2DXRVb6oX1Gz4OVa
u2AmOo/I66FnuNz1r1xrTCl1wb0HtG8NYbfwgQ6J/Kj7HNlmkQR4LkoIG4XpAH3MNG0yaUdq0POB
trPFu4qgWj4cmnTURzeVZIsXO0O3IB74lZzLNYMh+lcQVabiWDPPkS6tTiuInM+ckrMqyVovWYry
y9A68RBsI3cdXjN8aDCNWIO6TLcvHfdFFHZUCMkWm29zOSIGgzO9vb7OPv35sEd6uvhAoqIRwbdr
qficzyfegwO4nAYFHiKDwZngDrM+nMqncgkAv0u7Y1swQiXH4hK+WnUCbA9SMH80AQtlgx31HdF9
sANrk+UZhSLxggkWxOZMrpnvOMBsWexDl0DyPX+9KiRXNvHKtJgR36gN15B1vatTUD7ndwAjS6tG
njXgEJgLirOTcVWP16rP4f+azdD3t6AWj41UeduFwirsChhD9fpgjn9+qRf3vc5ctR3PwA/thinV
ubRP6AAoTKieGRQ0zvWXw4jxbK9vxolkDnMqhh0JJoU3tReErEmAtW5pgpQAUp526gjoTn5BvZZg
TiqsEc9z9q/c0uRdGhW4fNnlfaVB8fxBIlwJTLqty4p+C+ZptVlZCCj+nxqglzMwq7O3uk/9tc6i
vGU4zr2G8dD6PHBmmuXQHEq7BVeY5tfKnDxbqTmLzWc0kaGAiIWbP65fLt21aAiw7c7BaAG5lVxS
GZA2Rvo82musYbEL1RimSmye/yx3JpDpDvkVZ+5Vma0OCD5YbJxPkW9JcxTWdRVO3BmioVHbADFF
J/wUf5AIeAA0nlBr/EgVGoCOghjhlLQK1GJOvJlza1mKQ6477SvbInqKBxu+XuEGPEqbAVUaWGPS
AtywIXILuoJ1G4h6dKz3bX6CXf5LTpWnWCg/tYsGJEcWeiVNLAZeb6AdUrTcnbclKQnMTB+e3pNV
ol74ulOQWaaTO9YfXiRpMCEJ4cw2znQIcwp+cyE8DYPXGTsjs7WsJUH+ggNpxGcdH2OQwAV3Zy9x
FP+H0dE4hbpmU/CfIIyn1miFjpR8MIAAucyUVMiqQq6E8q8/3XGcjsWWcxuNYO3ALUfi758ZvyDM
hhJWPa1xOabRmY2nzBrQDrLieDYx/xspsGsoTt5I8DKqd6P/R28oiBPkF15o5wyL+on5wte/Un3q
0S23VWVw0riBkZDFrik/FygODXOpmAPSN2mAB+TqebpxYwoOCYEGaeXUf5udPCdKKbXACLENFSBY
BbEOWFseQRlxt3X5NA76IHoAfHvJ+Q111PK5LuteRWQPxuGhvTJb2JXzDeuXg7vEHOz+IcxE4la+
LA375RqBRStIaTaz5zQNytDG6FR5czNhGw1KsGdpLNsktlAEg9utpQoUQpjNxmKfu5WEHNWWlRGH
o27a3+6cx/BzX6wxWR8FA6h3xTuuE9XUgeZQ+JbYbIMdgSsU69O2MjzcS16pN6ySRSTRyb3ZEt1R
9J7kRCzVhNEIbOO1mTB/0E4mIjLq+Llbeg6p4ix7yQenxNNUY1aCwnl/X6wUhJp9TsDzLRDqHrHR
Lm93mnhCxPPo62hym8KSPKojKkTXjb3/ktJSp5DJffJJZdcyOZ7zTYa3no8N6imlXybZqZCt4Qps
Z/gsxOaSdEZJIFr62HLIEa6vQNHaZtdXoI7LZXkTvW3eDR26f0WmVEb4v20+JIQ75gHoOQMEsLQ1
37xSmzgVQCZ7kFurOOyXtlk61DTYX4uaEJZ6UGx0/82fc9wEPmdYuMCMlwRZNnQ6+FrG0tbkoGyx
ZKwggMfG/vxEd3IabNF1S9D2Qh40zVmFxHjaVT1ENqRfRiH0vzE6mkc9KwGfwNh30P/tsp56X2Tm
2EPXqSGmraO3JTnZklKMAhqU354b5pa593jsP2WEhYqHM3yVZCiFggFXbU8ni8Qst2dWhAu6JMcP
SrqhVO2QJjUoFRgDTPQLeFXwQGBhWkzPIgLMCgj3dxuRjXAsQObIzM//4cccNB0dGmBU/35131Pj
3R6N7JDft+satYVj9ZXp9Op8ZAQ6shOW+scdAmi3Tp/wfLmLuuDFiC/6BwQ5eHh8sVPCfhKcKQC4
4j44OCXT/h0nAWxbe9CDjCqyDypaOe45mBWW7BkmGUcIwbYTwaKwIGhjUWlEbdrveo5quINXkoYg
h4UNcxLyZqZR++NnjNmFJL8HkbWIz2cVbqxPqoqPxWxpaGGsWKMDVbW0CNRoE06ZXAra1q018WH6
hBkYcFOFSuVB+700oRG6SCvQbeAVN3nUCbJ6RgO4UYr5Li/M6KUynDykZ+f3+kBLRufw3LzzxPlB
E5/qQJaih+l+Lx/Id5cV8eUehYeNngWDhqCqHO6PmyJk+XeHYW7WpYsR+9f0j751TUXJKiUdukRK
qsptSG57oLIzgvlKDXl7zvV9q1qSuWQ1vIpOkHdq3BvTMRR3niuLJYXSo4qTEvj9HSjxatHl6flA
08rqoyE0YtiK1EBpgtVhAoR59NfTGKcnCP5jnnucWJITXUiPegfHTLgVP1foDL/TAnM6ExSGBnWx
4d48SLlr/tY/qov3EKMTXSyX5k3+GJMoFE0HiMbg3/UQSmRnEDsNOcbuhWuQBETcMNqqZQtZn61z
TbsgHI2iNNvMPZg9TgpBDsBQt/wtdw4kqhMOSghQ6qWqdgspYy37NuifHlIFCc/iKyltzdR78zSq
r5RwUkaovjqSU7xbte4sTNuJ3mrlQg18mUEgdo7xLYP9R+R7CplNgwEu6rAEV4OLHUmRiwKTYzd6
9fBt31R1Ood/u28zrVkhehWv1XhtJ58GcCSXnwi/TNcarMz50lYzwJIfR22Qz/OeQZyBb/aI+hrs
mQdoJb8rycdSCm3Rw6OggibIBGT5O9vG21/i7vrLZ4v+YJrIRFEgfE+sLPe9O0gIOt4qDeogkJat
SRf2v6joDUMrfEIfoFFTDWRBZUCsJ11fv8+SztJ50mnYg4CPhcSD/L4ogRMY8/GZBM08VfVPHhpt
A2Vlplkidq4oiu8VptxLZ6oe9s1MWWx9OBxNboewYN+2SKe2KM1wFPV0Yxq8EJ0/s9HXRH45n9hx
S4oddW2UJ1WvQq6hScJl8KZWB/jWLb8u9ZY4lrjLvAtODIr7RdxqoJpgU8OR2wjOaLRfQlU6uCW9
NqFSRoEA1uvsHPpEVAdVrtSXA+LBDGD86dl2cH9smHsQ6j9HRktTitdiECkDWTDWSHDfEbQYBaI3
eTPUBRNLtuIPR+mQuI6gTfKZv8xPswBbVjPhmGQa9FoHMAefI8gnsfLqKsOEZ7YHj2fZ5o/r0cim
92+o6Zk00H2tl5Fr8owTrDHPL8ZuXZAHNqA51FTfe5aB+T5vxqngMmoPL23mDq/OROjE8BkH+DZX
2Yy9bca5f7qd14scPT3ryhDTp5+BmMyooYTs41JRveA/En0ENfsZixGOyb2ag6fE5EffGN/eCjnY
1mmcfAoigR+KV31xDeBUBsQ571JEDMETjFH4LCXs3pA7TAObEP6SrhDdRHuObI7BMMSvZU2Dfiek
uugONzp3jwcT/k3LUowm2nNgjPo79yJZHGR3l265yogjzoUxp2MRuUGmjd6H6xQohvzuMsDYORH9
m5k8aEkW745D//cnbF+BYeu3waPV3/Yjqga4pI0zjNtpm4LmgAGiwKAHVMmXatWJ/62fjtcyPzvE
9vjmcSsm5Ka/L5EPMSi8jxzeskYyCewmWLa9l/Kqc/oaQwb+b8BmFGwzC8wJbEXXSbxEXIQO1h6l
8YiT76B6JFQOc5BrhsHJgA79ir5OvlaRu1ntYgfqW9BwspkaUcWIB7J2fygsNyRmFE7w5TVYBbY9
uuWs8ygERqxCSqn6TuksbAxhKVFuLYOCzsFiqSB3S86sOWD2wj00KC5DYIw06MJSepFa0NmGEEoZ
06lkPPvjbwYGw29Fnr5zicTMB4SooCzbmmH33UODa5zzKS01ZqKhoyc2Cqnji7wIw0uoMj0c02ot
0K4g5z1x/WFveWgWcPKtgPdb9CDMpPYoIIRdXt9DFxjUT0Wb4vuo8XLnmTCVPaAL8vueqq6hwntK
tCLrdQeAZpjOW6iUr2aklTUTeoIdz0xo0ZFel+we9gXeTrQaxp/00M8fcP2WSFcRzkcbv14oVHUs
8MxmVXaYoD3HLOAdA/hA+fw6q635fNMHtqMCDsRXYCSUVuCuFRmp1H/xqf+ACEH+EyL+Wl8N9PeP
Z26twkVJnjXSNGWluj4TflUUPPAgyFlVY7uNxM1ejv//KX4ELjR5YsTaVtQROFNzlmZHUnQWQ2Tx
4/r2FPzpRR2JUsK2E6dLrbdw8QCXEPAqhiuyKCLL8RCMvFSD6AEJ/7RSL4hZy2qnniez1m9IpMPv
L3xZ//eGtge4iPGDBD5rrafxT/YkcS4eeO7uYoExueyRmx+Beds047mOnYKdxrJLgU6RhD7juYgf
ap7f2gf9avbWnDyl4N2JU3a0a41BdmGjE04P2T6xYPWq//hMfQfXlVopGfzNIcEyM9QG9QVi8Raa
/DM93q+fHyKViZsKkVdzMIpgSvTq0CREHa2q6NSRD0Q5dqWYOlDWznWmw26fUhezJBNiiG9D9dr+
r141/u2u1tSZBVSWXC5Q0wiOFdvpDDf0fBbzSgU+P29d/U0bPXfK8jW0NjlMuQSp+uc5vdWLR0MK
30yKlO2hDrRwkAkCXAjhc0Gb0nxB6wk+Fsr47b6a1ticyrI7z8opCdRcRMNMwwhzqqAHo7ssygdI
jAalPzz147A9tLgusBahhX8kebSKUoZHF9VuyjU4ls3o+WNiPDrsnFPyHJWhvynCMgkeQ8MCR97n
NciZ2i0eKD/Ma3UN30wSd/zogdGVFB9efLV39Go6YiB/6kJRhscbXaLPY4BfGgplbXfsw3rv6jG6
5/IupZeqt8Q3KhfllNjCFuCouIgneAj1hviLH3fTaOuMPeMWP+LsMDoQ89s20JwSnB5+jwFgXpAX
nCcDZ4S68enAT8cdWtkbXhejaWj6qTVzzHWW+Zy6IMjerT9XP+HrDikt4HseDwvChM5BBv1WE2lY
02w8foyNZK71uevdDSBT1mzi+dgIp6rb01yJemGJnrP2mJKPFW91QvjGpd5/Zzc3n881bYKqZMMs
vAuOGoaY/b5HpFwn2DNAp0uH6sRVewvD5A4XnnO+OtInWl7RKWfsb9MGUtj17fvYHFbdouWftGuE
AH52eI4YuxqwNh/DehDxyEoVbGN+T4kYpP1fk7Byd4ldGra4Ehgq/L+G1yCW2yYXUIOlAVaR5oe3
BCSqivTHcslckfPplvRDUJBaiFbh4TvQWRyuVcqcn6TB0lDkDid7C/vn13wATQEYRBpWc3r+tI0n
Wnf17Bw/oWZ3eCxg9NhrTlWrywCTn9uV75IwWbLj96s8X4A4hNR72r1/tPGCFbqfDLKX87C0zOXX
CPO2FLctrssWmRNe7dTSXdsQ8jcRwZLOwu72VXDLFW9zBfZaJrIVuIYVgp6I1CZ/KqyCIMi8Xa+Y
KPtrrHVCZoy0OGycJatJY3JDSrl7diDj+DT9tLmZG835oMeqX4crzTxpASsLStu4UwqBPfM9vIb0
AL4iNgGo0Tce3ea1l5I/K3o6zigwDE3ViQBbtqDHNRCIoQyFFmXsxWC6rOcVATbGDul1sGcD8kMG
aLXmsFItKh3EAD1etu3AeFF7uKC4LH4mIe46xu3Ajh45RbwuHF3G7RVCrzkBllxBAT0+GtLTsop0
oVqo63KzNJW13SsstsvQn1GrcUc0fwIhaZlSenwGoZ3UpvjgZdAvDLZ6mEHYn6G/nhjcsO+ccGUK
BCiBdk9/7H9kEs+hB7ByCCjjVoWzEhhmrq7oh69GTfSXm0Nd+FVMK/xY5898ueQ14RAIPK7ROE6m
P2M5w5enRPBRgTz1+pa1tZak0jpaZ4+iKQRWr2z8lR5PyNbch6DKYkKbVKKtnXVZGEts0t2Ah1wd
oDK0PyPHVbgr4UeYncgAoZu9ouBQtM0xV1/E5NesQluQthFn4s0u8JvHCScDDiuiT940d2frk9xz
gLXZRy3241R4BhilpPtGHLbGNjYJp/aV+fvrD89G4g77/KQxtz7RglAOOB4zm6CKKNeFGkU2leSl
r8zXwKurVUiDpCIruejii/RGo4zRy7b0srGnR1ZqAdO2N/VjT/WGLLqGxULuGhhj1F0/6IuSDr6Y
35mUGDQKVJW5mrvcWLOAht6FbCFqp4uO4KZwilxpNmdSDdkDYk9XGLJRKh+WtRBE40yWKVZdF56f
v/6T0ZT3bsVC75B40f9LwVYVPBSsqc/xFTcVexqMKihVxMUNfp0bdYfVtIXJsO++fY7Y1wvYFGV8
dcjERrWTb/9nXxG+E/gUgjjZDTiv1HkdIcl85ExE6q/Zk7pdJBpjTabUSrwk7pOWGCCWTlIW8QsF
MBVCtvDFZ+bpLuKc4ElYgVpgQLqN0YBFnUneZfG+MdV+bia2TFS1Wcf74wYW7066az5bN+d4qVS0
Rd7YuOfAKoo/LZRkAahpHA/CXJq5kKCCC6G567VbmO7JX8pCkrXFwPlRIGcjOO2XwsakYq9G01ne
xM/bwL1zif4DqAqRucmnyBV3cQzFXWSNLio8xb2w+Sqzpw0ZsuJ/7HkhZ+OB6s+/+1sF2R/miBli
2k6ZBWr9nRrLKn0GK9wovYOIlkI/g1lF/+lj9DT57Vck0GquaAWC5TWuiMjtSLmK5BCJApqtyWdF
naXVuNhgLua1dJfJcgsUdiSMcAXR47dnlJ3/Ct+kw5QzteKiRuVCNrFCEE5FInQSdsXnZ6Ztzo17
5deMHR4ulR3bRsMq7L1Ye4uPi4/hIQMDUY+DphBX9dRDykRRaXhQEMITaspKmgb9c2prK6WZPXNX
N2OJMBq9uS5Ui/VgDSzStODS+fT1iBQF4ktWLcQ6vmVUE74G72grJwrseL2Yk2iDETupDDjqt7bF
QixjdFoHd08LrtWXs8oEePetBZ6diAJYVSlcNMFcpyY2IZLyjkjr+g16JnSsYAVKYNhwIOmLWUh8
y7Lj4lCL9lUmT1Z5fDNuRNerHDMzTaDgs53Lg028w/8lm0WaoEGFrD/6ZeTMTW4ocwbTSzjOZbvp
30hYQ0By2xTEwfQPMZWwDTgruMgvITb/iUlydS+/iKJgzL7asOpqeub4Scsqlrgxa4SO8OlN27Ay
ErhB6otQKKl/X9M24CNtWL0cyHwrVrJHIJPo9OUasFxr0dM6XplET8Pwrx1+ekGN7/Psu053u0A6
8SDM31N3OTOO8E2F/uRIG3idZa/ETxTsYRDWApWgtupx/Nz5N+QbFFS74V7QhSQh34fOhzhCYkUE
OveVZbigXq8sRP/uWLCntY15thHriDB4dsrRScDZHQxK/P3Z1oCJEfjLQ3+IcufxVX0pDMRhoyNX
ix00ynrSUy3+agBuYqS2rXwFT0rz9+yrb42PG9VxispTeinUiQfBYj+aochNqIhER7WS5Qc3YD4w
ljXd2CyxEdqPJzDZ5KkaFPRobHI/2AEyUB+Mdxn7MHBLniFevDe3mM2iBufEoIi7vwJut0xLChfo
WpjvNVmCvf0pG7vWAVI6hMAOZBwJrOO43XNbO9GQlzRw3CxIGA17akRCKq4Q+611svM2JjxCCWLT
Uwbd+ZPWKZiEiJwZhQF/ujEFIqbYWY5GM/O7NAe5ofuUGkJGIDvdwEla3cB7RhShqkqwQO2O5UX6
+8cGe/ay7yEGSH3Ou5yEiHSjrpKELzp9fvFtF3/KJh85Az2oV8RW7+Q63Q2rRz/5sb0eoTFM5vcu
u6BUWFHErpEU5mDprOeBElpylb3yHELLcLqvDrQqY9U6ClACnvwKS8CbWhhnnsaqbB1pyd8hNd/z
ykj7U68FgsZ0WptVWf0vbCJ5pyte5AgFsSppGcLt9g1566mvzdSR/CLnvW+HYfQwkXgiC2vZsLRj
AiguEi/YFMliK8YINiD8+inRNKkBGgA7oAwm7xJGn0uA9aupBI0cRxOx+rm3RMJHk7Ej+8mdH4d5
lvkYT05Nbl9Exr9Hur+++seGrQ7ZjYnP+tJgy3OK1i12FEVCOa+GbKpufeG6q2M6ADV3PRSJgESY
hxLatesHIckNnZsAkecnlWA8uqPie9OXBm8MvgU9fu9jmt/tTKcMXPyU5afQ2pYNOovXF9AhdWpK
o0tOMOgrLAatQUCiwryl7FZKAa/QpBQam3t1ha9eTlqdQFr5rzlZUgWSIje44df8kL3z3uHZqXxB
ulUwIdn3uWhl6Ezn4/my+Xmp37NZdjk9k1zoemEdeyzsbrBXGC/8BG9jhA9oJEfgPvh/qFyik0Jc
S6zclQaZMziqlHN6EyJ+RZbFpo2nGrF4AImZ+PxbV+xDrsl64zAI614dOpOts8RsWj0ZNicnmLQj
tRYJOgn6cR1a6ai29SYc+rkrk0j4XKusLEP9zcX/zUhhnoaG8cAn+Nux6zfKUmhWh3LwTRfhaoK9
XJAFr3D0iK4xtQdtYyAQqdHM9OEfbJY25HMuWH2TA0sg+mjwz7aRLDBZYlflqNdWCgrcjnADHlkd
W+Bk7OI7lhhAhnFAEMyyHOfs2HkuEosd08OuWoARtG+nOMK4zwJZYTr+lCpYRg2mqOsqMRuPF2ou
iN6ePdA1q4Zum0PS0UISS7cp4b1QJF1dBM7HniKgPqL5FetI9wKBAFc4uo3h1Y2wKgepLBdqzkvl
niZYig85+fV4BItBFrbPXbDEmHgv/m7IdPm7HQLd/heEMqTuBMN0/Kld1lf4UXVEmmlpUUDoHCe3
G7KkwFa6BNXgu/V5nWB79rOWTrvBWoqM7SLixDGjSHdZpNxg11ZuGGc7WG353vZzaEvZOwK4vY3p
9rMZfJdhrtJSnL75F605CC7wdz1Q+aTFTICg2dz8v+WtcIHcm8VUnSlZaHzvPRcHfxhHwtwZJPnq
158hkm2H7TFcM9djwZE4rsHT+8qMFaLS5YbXk3iBS12CHaaNV0Bsf90af3YsMnnOK6j1uj+/GphY
qXATfb51sJ6IbyL6zD5TLWNcLIi/imyY0zlkhd57XUvmE5s9asYN4xCz3Qx/Y5W0oAMQd7hA+cB6
DKTu9CGs3OpZ1ooBNGyhS8YzfwDsY3VbjVv/LHiZ1oEm+lcLBvja8kQr9yeI/Q5QdYtG/T+YbtcJ
554/HV5960iEiUX/6lpux0TkX6SRTh0C1rVdD1R9S5GegeDIY+0/fKyKuvfIljWemlGFVOa+uBKY
+itaJBaMYkTonbc3qYvJhRZtFKUl7dSUzqeTJ3wNizZ2tyFSkKzjG2SEOYsz6it45zSAQAhsWTVN
gMvNqarR7tNiiMQqZsWTOrPftr5VEW6qO9zSpjTs1PfdMnaykSxOHfREWzYQf9Yxw05K7ZU/q+j4
atpPIRUl67TVGZGCWlu+WOk+TrTdpf3apPIysPY5pcNMZkCdIp4vHWzbi76bb/Dw5DaRVASefsNR
oU+vp7RsVwss3NRvwXQWMukAU/73ULOY3PXBBqjJSCYfq1GZG7yD5CtnEseDqy/zdwcFjZ2FZfhb
l7rssLyVxJOg7mUV7V2rS5oyVEx62nwG09q7GaOBTt19UuCwh6lBRg76wIkz4Ch8AzPyK+IGbEdY
VG4yAKlbWEpBG+9XlKwXHOQUJmLKjCCIQkREWqzEV//6sSE98b+8PDKFi3QKHwHR87XJzuMuI2p5
eOzXt08ei9TCQqLbZjIfND9zy5Nr/d6JjLK1BR9tn4C5a2p6RDUJSv4l9jhozF/+j/KJrXwFwupm
cJKcHerpn9+uQUTP/mznQBFHpMx8t5Aioc0iy2fkK5DE1CUrGPCfXPn7sd3htXHvSQcc1Yp3ftsv
+UogFcoQxrdx7IeoN5c+gD23GinxqR56OSouaT2PE4MnaP1kr4VkNRXDDFofANGv+Xcz0eb0WbPg
hN36wleFGQMF9jMg2IwG5JbMUcCoSWR0jy3NRe06EwJJTGGDdklNfMwxGBsslaIvfdlVDhW9/4py
2b1SFZgVNrBqzwxnhYTQFwP5IiFm6fkMRrUxrqZMDm5PXzRXn6LOlb+UhIgG8q0uPJHUExPBB7xS
PmukWZj10mVBJBH3hIrkRWgIN/cI1+JeEMjS1znEG+9dEWN1qDYz+8hQbmh9+73GXHfLYTs3eKCP
mhWl2C6div7zyC07n3pHdTyPBWJFLa8CY++E6kiM/QCqIPCm4ZxG1gUI6X6MkOArRY2pFixovpPF
oVtMJIrgCe4NpDJymyK/BRKocQXhu2H58EWZSBL7KvC3pwKXCOlIq+QpPt4LGxkwU8FjwW+IADSv
SRZNec/ECp8Svv/JXHEiwkKJz5nwDKRsOWCswNu6LYiaWO4WBEx99AEXWCtsEGAH8frbU0DdRRLj
D50UvoxkrAYZ9nWLQ2LVh2iL8tSfKh5ifbZX7VJCcsYyUKtav/Cy708GtJq6JSbL09XjAnmqcdRo
QcrhgqI0Acz3c/DD6atgcG4BL5EkZp85kfJgBNAlx+nbAQkW/hJIC+D+C3mAqt30zhnx5ebn162Q
JX5ywUCzTaIkmSq49T88fhCzE5AncZsWdlmuMkkp3UybUwU4fRIkWzaLK01n4z9MbTH5lKUMdrCq
a4Leiyx8VKVoe80wPk4eaO544GoqtzG7N56kd7SODfHoiH8KsvZ/fKW40BEwrUoJYMqApqjELqVs
LTdLxlM35ZIbQtP3YYTPQmxHK4HkXbJWBH0v4VIaaVKYSQWKhqCXYYC7Bs7KGKeN8TBYqjT5vMD7
RHaFGrIMSCrW9C6PrGyouCkeqEmrWB6jLSuW6L9gYnLMnXuIMYhJ8PKFYmaKLH/0dPtvAkOygZeR
Gq7M20oYB+dIqHuzsXElLpK8o1MTQmKFegdcBjRci8Ys9aS3iLEeHp1Ige8Orkfhw19/StF0xb34
xYucC9ZgElNfx13fhdHRitF3kjt+Kq99UDIT/evY9HDSMTxePAMp4vGg46eFHaI90/pmcXDEsQC6
1JKiXPMTIpinTuWF7rZB/afGQCn833ScpTiJj6VSF2ll+w1AhIJ5DMZJP8QOcDLpV7N2VQA3mLUh
eX6mphHTijOWUEzN/QKkn5x9CMEQ7mpNwiuQAYY8pSx/PZSkgnOKVVlL7wu5NqVef3gYYOJS2Nnn
rmzsUceFm1EBWv2atApq+zo+QNgw+/TFgyUn2SsEUqveDxIzNpXnrUuj+QjGxQb2TezwNXyZXiWY
7JRuXN/gA1p6e3c+CvMsGQBHUOGeKWbL5dOKdyl58OOwfu5Ke9xAJjTvKOMrwUVD91nE30fYsAUg
HPbIxrwKwhSk4MWQbfPXAVlH02hH7xpXgYLLHN6P+wtHUjRFQJ12vxgUlyfQzC9lypLl9IWoTxEQ
X9a7c0wcwAI7Y6yeRjL3BZc/FCxr/nElFBwy9mMO/UUSbMyzvJUYMTPHHrk0jQoShItBfgWAL+Fj
ckiIeZqUYzW62NHcxoHOf6VaaQg8zstpIlMh8Uauhvs2VjCwwCaO2jWUfx5yWtjJyKC5AkintpBa
wOLTAJbeE+34U5+YJ1cbfL4tfyQOsXZCI//6amk7j1yE4syicFIVUTdoV79pnyapGWMF5RGzE9z7
NWfxd6VgOp9yHTLFBUvFmro0E5F7t3P7TpDqyP1CV9GEj7mqP6Of/WwM9fqKe2SpRCZ2gdTJZAmK
Om7iPrUWHkqSA5AfImdKCq6nTXcNcMY6N9HihcrEnww2j1PYXA6B376C7Qw+t5Y00ik0ITbEUW2D
rKApVUPEzTFi40/7xJdtY9M5+K4vrl1X1p4o74KjZWhJL0hEdClamnxen9tr8ZKsfHUCGC61pilK
XN8q8QuHzJsSyEwvT/aN+3fLJGcGIAGmZ3JRJPpOm9mhAdrwXbcHvkwdyFKsy1dlnSecHJF7sdYh
jjaR3zdgU2spvmeubpxXXEjm/Vkc7FHP6HrgmmE7JjM5BA/b53rKTdW9xOwSPEnpAd7f2JXQwNsZ
ih50DnFV3diocA262XmullXJKPN3H2UnfHRRpqClhlKVueCMopcvfumYlAbOyQcrF7FeKoL6KL3K
wtkMyD6UWZ0I0srx7Kh0THrjvoOiqbUVQ+TkPABzSdHp+KIFj2BZKkKVIZKp/w4Dd0+ZWFyKfsHY
yNkEjK/3B2ZFzdttr/Dgupn4hj+wKkpK/YbXvP+kTIpj6qvGJv5pRaliSJ6pPb8pQFjC1in8gFVV
jmrGE1Bq7Saf40rQ9Kx2kqMLrbJobM01apRmYJSTdqe3wkhwILlQ+BwUrgaR8u05Du/iIXAF88hd
OJvEJIjrYZVPkBm+SGRBwXsyG8iupM3bQnsNHsAilGSRyp6IJR7GR42Vb41OQ597tJPH9chSWb8z
B3P2ctbxFXhbhjAcGyExgpvVBeChI0YQjnO1O5M6znW+DtpyAIK0/qMEZzh2yD1irGkURLitK3kV
KpdETzGpr8402qu+u7OEJs/erSboR8tsnCtLGpDysb36poulFDlFtMHK7gVvpCQ5FgcFujd7QOb4
hWmacDlUipWm271DcqdA+YuiI1Ab38s3nG4aG3OyYC2kQ5A3YZbw55TWBk7TwHxcvQFHQ8dILDPw
4VA5JpSCEzKlfd43+w3UXeEBX/oxCV49ugAiI4Y9jddUAnUs4clDIIAda486XkHyNGR4qdukBied
RLMIzz1dRVJiAtnDSv4mpJ5VbbL6h1sIFJIvS6hHi7jP9UulB3rRaDQAqQjnMA8e2kxNQ7I7Cr40
cUMZkyMgLoAWFddd0RCKL141K+l6kvZfhx3SGokhY9n9elSaPWPGtTYcrwLBLpCiA2nAd1DAqD8B
J21F2MHk4e07QKNI23C7zskslBLipM051vKIvE28PjD0nN2ZU5XX2/fktwReBXBdlVkJzIoxKfdq
4NCPMfDU1tI216KB41E7Ub9Sz40rX6d0HvWQajWMTEjts08eOiVi1AiUVuCsVAgR38+bAjhgU3nV
e3NmM0pcP7vw+4rRpSVcHRHbwcreKCjKWm7wxk9wn5+V+rMFLJ1THTmkE3DAsSzgACq1L8CvbPZ7
tWlsjY1e0hpRfuyTDOTed7pQhkCupOqsS2/DpO3ygezqeUkNi8kNuJiyilv9l3twc2At0dHp1+Tv
YGfSQwLdQLlNWNZwIgRQKgbIZGzdAOt9O2BREnnIEifXj3NZeE4CphcpPDjAi2+643+cJMtSx4WU
FKevj7evYrBtZJ+Bz+j0/hNhHR3D8OXPBZAfV8tv4kq5M6xwuuJrlbij/iETXFlFp+GuUiCzA1Uq
fiyroclwaWVGf/V+2zFLiJPRIH4PLRf2i2mgBM7jG3LzGWTsftyuvXhZFN3pjFDx6gEYuINQvGeG
cGDKGHLW9ejb5jxWwbnups8xBvcj6uKO3Eh1bJ5yHqyBfT22ynjb6Qhx2fWm2nUlv5ZovP9AB2L2
mLlBkPoT/k1PiTn9mutHBLrLAk0SoGh/B7JPWWzgHGtCzViWSWIcYYkmsDPNgM0nR/OJRza9vQd7
eGco+320QEi3IBqPGzjKcB9URpdlOBVqQOv1uWp8QBNaQKSEsGJb55yPGCc+pcU73iK52SxMwdAE
+nhWf5jtvdAFt8AuV3O7bbG8LlE79VytQ1dsrzLnKeRWs6C1fXSMSiNDHzp7p4vJAVK4AARn1Gsv
VxnBpQoUgnjKudbbcAkjvmROJJy19spaW+FRfaoRIqgLlEEWAWaMjiF/r7ElKni7dT0qnlGd8zqu
43BK54pQ08OOGe4nRuXA9jPYl9VHUhsS2XBvLn28O099btL83jbYH37PphpESLYdmzGDqRypE2EK
biqad7FsiKqvZVqpZmizuvtrkpUk/OxrlGCJLMgLqE+jn2sKAV+1w5kHgJLOuF2WHdCkTOBKh1c+
g/aeNBxEXM0Ua4LOJELtHp7ygeK5I0lJXc9yGvZLLm+yGEV7S43L0FHVXp16PmP5uyPBCp6yhaaK
ZoJGrhPDSLKytrcDIKchVSZpRV4qJL3b0tGjdW3RfwKXUSFQop1cf0TnWAEWQVGGZHEaZsnRLIif
AE4sNzlxCejjmXsZhkaT0g2XKa/d2vdvmyjYYSpFG+fxfkSSNInuDjtltyE0xmh1oSNhYS7zVZiz
OSAO+MfqKaUlz+bXODwrORwN4cC/V4iu+ntHLuftJWqeL1gGJmjHy5sg7I2HeVwHa4qrSxgCBW78
tAdf8cuyVKqbGFBILUPcVVVyctr0XKBiZ+o2JrZOW4NUyqo3hULCDjIVOLWRUqTgok5W/JPDK36Q
ceEKnkhqqzFAIcKlF6WVZUEDy+NYK2cBKZuaQbok7LomMz/OIcdN0+Ji+t65Xe/SsrV12CyAgoVl
PE+DLdg/maiz/5V2iReHOeNMFLtSMHaJ7btPxrtaO9qMUihGjsaCf1DeQ/BnBPGKGXG/cIf0NxDu
MC5HcSW8J9mnYlwLR+OPaAKkS15mrSQtRhCg6dnvcIhcndVtEwzCchC8AkyKnKJjX0wHy7kK2yqs
RVkZtSfxGEP2IHa2NG3SkhlbyoYuaXWGRtStS75GsgP8WVXANXWI4+9IpJD+NpT9PNPLL/XQkJTS
VG4pqUuD7auPe3GIbROn8eVF0IT0yyWvNuddE6g7BUGmGrOASCte45Yrh6ovQPqWrqg/1o4SMQ0Q
DAmI9UC3oeWzuHXTrH3t5WsdyBbGNwayzRMxxhFu9/zFHs/hkLacuFZeto3o6DxZFaG0s78cm2YW
BbwQ/T5RUj3UMZ9wGiCTOirowU2gMVA1TbsLhEufjfbLrjol/BUTD6m3Lfqole6UDqkJz68OG/q1
PSYnUE5hnLV06K8HBEoPpP+n42Hwbo1OzgkuZe3OdX9PLsBQHFYREyhOg46yiW9VTE/YlODR49Ru
sfO0Qwp2GHjL7W4PwvYjmHLICzc58UBWgqGtFIxOVzSyMoOaczZCivGp+FNb6pSfLU8wiXddEv6a
11iTowIQbtgQaNH6HATK1Jn/be/Uh4TAaECI1kUBcKvsXN0SdJwO+bCSW6tjLJ3yf7UnY2fu8OG+
rvKUyvGzHIr5imSCIXVPbMZ8nChfbARo3DTyhUoVRRlJk2x/wpsk4zAkDA9kctbdrlIVZTYViXiR
D8As+POS5XLh8qH2ZJsI6uSXK5w++QrQEXogiYulLH57J9liAjIqftZR8Zl4YhD3KY9r2ilZ1XQI
Ia3TPRAGYzwJKQGptcMv0tbz/xS3HAEdMobbmnHD7vn57mmauz8S4PZeRm9N/X5lSE42OKfNQGFY
TL5ZBtre2kp4wspVs3HQ64nP+vvY5Ou8rbQIExBsZFHuQzGH1VS0gWLKDU7LECyzxL4wD7solQvn
d6hucU+gelu9gveZR4y/OFuQXLqeaRyVo6bzLMY0nsFZCNl4nvovoEZi33nQqICfGLQXinGdNiQ+
2zuNfjJT6vfyA0DOetKLSk+E8JwgiTmFaDCSKCWymRMPAe0RFf60rRUEo/M2Ixkl9NNaTVQ+qckv
2NjEKSA70cL1agSl16NRwKi4v6rqp1YGTUczI/IIBvutxQ97EucWRR/zaC8004H7R8rYdcjHvfNz
OCsUJVzOUoaSV8bwjkjIGsJ7krRFcWJUTrcr+6Sd0f6eSGJlhmB7Ft5GB35jTef0p7oIW/pnHgiJ
O3kksMb0IOI4P27PJo8b0NSOwBe7nKAbzkJ+nYUnGT9ikrV+i1rcTlvNYoSJqeAxCDp2khU6xopa
r0whFtVdeqRT02iYcoNr7mqjJfhcDLng1EEke3XhYRXRxcKwrgMRGpc31AVuJprhqpQzSXqAno7Y
EfGKAaujusJrb6ZSXUONlvtMavjMsZdhGrjH09X1SP8fmRDDbF9842U1VP5rb1dVIDUEgDNxqOd0
JWg88ymlBHR81DLm2A8MbThSHfkNtu4BsiSvZDaiuvFm3eJ+3T9CbMCYRsicjqbxA1iDiaqArj/G
lS+kIFra72Zk7R/w2E41Nk7SuPZlFRkzaZaPW8moilq2zLKuH9OF9l9jVBwPvEXs4yNwwy7fzDDk
Q+1t3lar6Uo3uTr5Nxb0tmJ4MDC+r2Q4yMcb0GZEQnH303hetEI9k7eFYKDjv8kUABQofwJIyk9C
Y96rkvyZ/P++UwE6Aw0LtumtdcDiv69n6OAzfujn1PhNH95IslETAxdAxjK+VXf1mCqdibiOAxYk
f8wDSiFk3z+Q8ktcTOs5IZkC/ZSIMFYi8qDI8WrIfmdpfj+9EBhVEF7EX3uloDkCdBlrOQWoXANF
6dYOG2VFu+pVsTk6tG56HE4tfJ65lCqO/x6gYdUth9jR2+srCGBMGK+QHJ/Lxo+ET8g9NFWa81sJ
DeUajf/ydFCPQ09d3ClWsMHmeFWZDygx3WhlihzNLu7HnaULKsi0JqCKTze9fsrEoMlCeq8bDzex
WjofWnAQFj5SjbcKNRfnW2rcS1eqz/SAqwNIp7xBBvDXhdSFaf9hbBn7im7xKgKlxmSkFmkpG2zV
Q9QOTa5KAHnbVbJshek/brb0BhCIv0Ef0RJH8LO/t6aKza8WYEWvIBpi6ksiWHw4lp6pFMpr/pT7
Z5pXfUka05BBRXE9gtoduRa14+SfQDyaN/+vOe6CsXhzE2ijCNbVcCEOVfC7PTDWOB63q5pZXYAr
/9YJDYXgt3wfWpMT41mCg5z7BScB8CyxLrH5RT5r/Uk7tzWxVy3L5WopDt7zUaHFSJV8Wzm8+UtK
NNqKkcBD0imMvfXfS6R9Chq9w9om4GdZZhY3KpJVtYigTz7acSMOgDySSnH3uulsi7oBhmzGyVZy
xv57vZQdJm9qGVymIYBxOqHXi8IcX/FC30+9hZuHPlnCzVCWA0lfRWPlQxi68eLLPJdRXU9Y9m7C
FLOHeejd3kRrdycJN+LeMud6doyX9gnsAk4Pv0yLcxCiB4Bsa7hX7oOynAPxfZ5pch1l37bEJISK
Q8gtZ3DlY7WkZH0uZXCxFGHmTCx3rX2OilgZ3XUr56QWgWH0ITezkDAHR8aEnsTrSEXhCrYZJPQ0
m/LCpLtjXo+3S742aLoaA+OhFdgs+HPdpAF+XPGxLQkqHQkQR6R9DwT82ujifuBywHdHr7dpByAR
6uIf5nuYr7NJggEZtk8MHn81/5VVhqu0fA+2o61/wPIGoRN7c8f5DAiLTs5POI1dfXxBSwHjscjG
oQ1E2RM6bLgBGNeq7XmVG75dszxrQ1POGnNzI2s2nAGqmEiFtCFJ3e751BIWPDDTKwl144VIvdoW
soKBMJr2PQCg7ZTXh+z8HlbsDoejAPFLhZDr2rY8oBIsLV5hZpTawPRU45tjIJnZqDRRExGiWqfh
L0LzRo2HwMvIB5SW2IbjE1y32EW3Lp+weuvGgUOBa7X1foehyz+kNDT2CApPsizMdg42zZ+Dl3cx
QtnGRmIcKCiIaOU2tKELxV5AY3IJqeh5auYB4RAH3AGHDheGSS7Pk2lTDVujn+E+sMtXplZ5PACk
W29EqWgH5LhXGA2exhypS0L9va7vp7qvf88veqZzdlXcoR2r8oTcWSjb9iZZCgEJn8y/02s86HTk
WH3ZDiOnmcR3lmSuyb3ehjbxiizFCT6glNpZbEHo04vUV4DEh5ZayBN9Ik9CkmXJXR3FhYHaexrw
QafqT2bigxzEzrZsS9sqbD4WeqAxJMZ5JfuITQJk29WYBq9mn0Rj/3NiRdc+0NyYagpsK6K8kXAZ
WIPpOG5vO+8ogY5CgA/cJGb/AmPlOPLGwDs2TTMwTWqldWSV76mS8DwaDjmI1EPUXzD5xYc6lf5G
Q1hkVlV+9OW9DHa2DaeWObs4Jca+tRc+2ik7ON746MhVnFnj9g6yBNgRKXyv+JakjBkiPWOEuPSw
26ideMGQmGIbsMDw9OpYrzeu9J2fdx7ThKrmFb0xEg7IoykOJSFal8IcH3eo52ki4FoHhipVfUmQ
scqVwyE3URPlB6XnSFz6bpswwu5rYvmbRBj36uia1e5s6XLEcmQYjuBA5w0Gb6CiNaAMX6sIDcUD
kZttjNjaZTvXxQovMUbrzshxXyX6XMsVSI9EGNmoRKWCGlfLwWdwSM+OC1pEGQHOa1v2EIlYuDN9
hTjTJeXLX9rA+EZw2ByAmxOJVBA8hAOM74bmPU1d4aLANHcSVuwyKf2nX7VGApo7qqu2oWBW+Hqk
zyXI7oMAB38+pEx3MhI4IaF0gkbt7IkVUwuwiDT0goGJAeFjXSJdL5o0fc2r9VAc4Orc1O/VOCsv
uqFxsqxJgmpUv90cGAVaxhcarPX5gfLhu0xOlOu2s38IzQAi1SMTboe4QFOeKrABNIkBCLFuL+7o
Y4hRY/ZjOpblHkZXuYocdcmLJBFUFi/D15rBWS7jw3Gmq8qzYA52J8B0T6BN0pWVbKhVUuDr8ibS
RxxVt0cCTmMvkU2GurOK9yhfe+X5UxyuSypwfXwXs6QW6yxwKcmJSYfC+AByUNRlEO+GYZegMLbD
pVjLjrM5ZhKL6/sb90CyxwV0wj95aTQ7q1Nn4YVuZCCqjCENeHX/4lXCthWdMR043iZKIjW+ikVM
jZxxKXTeyITtrpXoNDs2sAOIJeJmR0X8OjCo93J8nL9299G8rA4QAbbaGRcloCuH2yPUAzVxX2/R
qt+ltbMOc5rY0f4olrPir1BIRirXUMAcAZKi38DRSEvZBu2/YOiOUFFjHXE9I6VTGLEzCIlImrAY
htA0y/Kn4nPLVSy7+YjHUi+OJEH5lQmzQTlP72Z05BIDdZif/ILcybG9u2liQW8z8Luwcg5dWlBd
qBYpbEaE97jcSMX77pCaPV2iqmVNkgZ6zI8BQIJt12M3dmp/5rJSLqgnXQTEXLG03P/VTacpAnLU
Ka8yH1LU72gtG/qETB1HAXMiuC88azhDi7FZoB/jelmADpCcTKrXhoHPCy/72ttjHs6dIP5WFWi9
qjEEL/YOCVv9ZV9CUZLKTbOan2wvOLfKC3ghrT8PvnF3VL7SQZJ47jCmzlB0aK/BpUSaEBHAtiqr
AJDQ4RXz/QaokhXb1CY1Hc+hMhmBzELnpnAjAQDMECbgeh4+9sNIGGUfOt/x0eBE+iqXLp+fzmK9
BMhEvZ/RPQoZDMuleboCuMcQiwNFDtVHUp8+/vDEtXQgLwjVlhfU4l5cuqXSv/8vJLCVgK/h606c
yyjLB9Q1xRA7BDPrXUTUQiWtEaOI5IR9m5q4Ho2r7j9XLBAVOPmP3CrvoD2GpvHVSKVjUb6DGdA/
0RSqugy5sSqm6KvAhvgVdViQF+sapntEMcMHizppF+W58c69pLPfGl/h+zFK9S2jDcES6FoatmEU
+A9mHAvK6m3cFaecOKGf82yayXOYe/S9Nf5xskD6TK9h02MRb+Hgf2srBLLXJ4OSfOUf74oHcZKz
5RAsggHg8cSIMPAyMLi1eutzopMBSxJmmGMLdnSs5AUMfSYRq4Xmlou+wRES25yByiCixDMa1Fv6
AI20IQQH2Tj75aVYwNQuVLMUznjLRCIVy2n3i996HQFsXpvj1dCgTBo8pEkrMrTihtBYC+X9qtPP
G3uaAULik5T+hAPU3w5hv6V3Se72Q49z4dV6aRfj7ixR2wShOHH31/42qi0UL0oDnSZET1snxhbZ
9JyZcollWD19cQf3p7/uBIv7BzYiSN5te/h1We1Fp93uO13GioUDTpzrCMP0E+lCSwZHNgxHdXkY
9+jQof+63dwZ/1z6ze7oWS336/iTBTcCKpm4dizVF5mX538Mlj54IpACAllo0tOsGPK/QQ8LXT/y
2Uaue2LDxcf7/yYeaqu7HJg1YuqotKS6akqbtFZ45e/cvD1JP5gkWjJgU26ovqgbayyU2M7VbJpo
Hnysm4H+qdBucljRojz8KUg9tU0QezmR/BHWjYzdpyZyq+vVcBcfPaSK+uqexOqWg3dKNWSazNLi
Zk9+m8Jdb4XGgZODRes2rs2IVkw3KeHYO16MWq8W4K8ezXoF5k1OFrCTcYhJf28AnK5N2IlU/1N0
nHy3ghpVO4FhasGYyVXOYbfbpZ1vQVjm/DjG29oUoYBsue9TWKaLwqCnRSXOpVS00JoIGYy478hX
UVYf34Bf5BAUdC/krcxhTXVs0/hq2laN+LXe8pgBYMZbE29Us7x0A4Sgfm/1ss9f/VgiWPpc8qpA
QjlCF8WtWy34ysNvE91cjoZ1UZ7KzLq4ReLOgNSzsbOb4GUrmJYe0eMk7jt6I7b6KGOQsjIasW6Y
/mUDuCDaGz3sTdWDfWU3uny3HLY6+GdKimKe8uVUPsiVyGzWnOT4syAV8m/xVmEfD+z91HrznQbT
KXY53uX1hec6tBaM1DtXZwEMHykS0qICesPVT0rMNbtOozE5Yo3TizP9ZOveKscMlsTgON1volIX
t481t2jPbDLKB3cmkv7E8XwCasTKmoNEd8CO8E5GW1hhc3mXNZun3i/dFAUoNFAZVmW3pN5b+L9j
pxSMiI6lF4RAUjC0IG/YYErmRFEXOJQrKRS3CwyvIhPmSoLz6kwiGt0ketNDZZ5ljErYSyr5+4eR
8wbe/cuXRdiuYgQHjHm6yhrFOPYej+jLQKy0fi82E3ZFgC2DQaVwjbnLUI7PneUD7njUh2bRCclk
RP+OiraqvHp3S4I/jDXTMgNb5LkwLr9hvZZnTaiYBUTlEO8b9RuBOvqYmMvzwkEyp/idSRLaKeaK
jdncMG7sn8WPewG+0i3WkyEMTmsW33IctwcH7bMfynyny7563ev2+FsxuET/c8DsZn1eYBwODzr8
lcrpMWJaTqvHXfNNUc2kNXK6IEzlyvBTHADMtQZbss2bChxJS28OJWZedpLpgVuhTSjz+g+YZgc3
gr68Y8c8xS31Cgr4TZVKI3dhxzCk5OZgc3ZTYsg467zpoLnhrTcZcE/z7DBRGtbg+pbwNdjrJRU6
AswyVPODYjEWbq0cuNTRX9/RNebxumM8A65CFAv08ynT/JuzLtWcS6d5yPLQ3E/OT/NKQP35cR6Z
cLvT5cfP9OsuVbfOymOAOY9o1szlwSswIuxlarWZPjVG6yqiO/5BzJilvIhG/vZQvmVh+vXmXlcC
5aOoNRlQU1fOvYI9BzjE6ljGDR6l9QyPeZZ33zXHtg+SkX/OsLwkTptursF+Oa52ZUXnY1G63qeu
n4c/QpPM1ch004dVSZpZyiLzaMBZyTmn3R4xA5q88XvnV/cbjkUOBUbfXCuWvyl004T/TiWVSvLm
VDDBCawIzT3B+mLU2BU1ZQ1I7DQQWQBzqMIxVIpKGSYNQmVjBfanUZkMHfbmiR0S+ML0D2xIrBnX
IKGol5YrIiXlKSOgWict1j4n1K88drUhojcfyruSv8YUB10SOk2HjqQh9mHrndZsf7QNo1oWMJCp
Y0KnyyH9fYBn8kKayw5equpTFOh1euWWX1Y+oFEm95lpqAvLKCk5DudYAvu+rLsmsHLLNZmhh4Nd
z23mDIzQVcW7r+3nUigKIW2VIpGjMcI/nUOK0348cEE+Ix2bixsAzplFPiOP3gHAmryEpw0D1oHd
h5netyxg4D73ZCDRc3RTMR6tA0ZPZF5LJOl9EQhxvDLUT+piRqyIkMjLQNvQWS29viAufOmzVCCh
HSzBvJa/sfCAvRn9einBC7eLQr3X9zFmdGa2kLTO2vpERs4ClMCfvcPcgQPEdMVYS2+GMuACHY2P
orz5hA+xg0+XKyCcgwMvVRH/RRXzd11ek8Ai97E+i3y1JMwS8sfwHW1IQ34jCkdQw5YWitjDKEPx
e/BZKQIdDasDbDU50BDah7doy3E2swhkr5aRS/AAc/k9tyepnbfz7DMEojOD8z2i3A3IkgqRnUL4
/G9tQ5VhIUUKCKmPX2oYYWDBfxxFUl3W/Wxiz8zCLSlySyiPuFbAXf6yYYgvi9gPhKQ+X/BuhisN
MNtvN71NBt+qMwmQlkwbsFIt+OBzi5nZXzPkXiWxRpQfTCiIQu9MK58JslCwO8U6/NEbvzg2SjBR
OcjS5HESvfFsRriLaxwMNno+vUPOkow/AL7iUxN0NvtmY6NjJ8YN3WhbiCeLgWn/l6HWyztgJGUp
QaAlsgu/WlZDJ4henCUq4ard2n8lA5/TSGljAl4M4lcxGHwCxqLe+Tid4Odp4HnPLCCjLpojSk+Q
9ZgAhgLWd0/BOE/PBD5ZnFzOKIA4pg0UpCU8fqBwuJnGI5HD7DC2Vae4gGLYpSTyZs/psGuEx1N1
fUA1e+4pbpFwVdXEZfNrzwkpkRnLK5PpKRljLvdx1OgsecsH5zWvOGTsgNZDrEWIc/+MhtS2qUFK
vWeA/E31QkfBS9ggxjAtkYouwuApPyRdhdo0Bz8H7Y+5k1hwElPDZpY71WWIVTbSnmAbnqvebgVW
zoIguee6Baa0rzG3IlFMjtpAwimOdqlA3dy0LLNyaiY+8pYgjXkVK2THJa2S3jUp26X8Q/tj8ofD
kK+bYYhZk0Nx6LiuUoo7kF2+Fz3edKzXMVSgnEnZECCB8j3w64ENEcyHDUSFgBtIaUdN1Wc+7FzU
tY8CtQLpuuuHQ5B6I5R5YP2rOH5jZaNC2SlX7z+hFyIdFS+eNVvOMYlXBS7hrIc9ZuhUAv8Z9kgg
18rpRnaS0OvJx9B2hqAOkb+dkBpC7Cr2X32QxeH9U/Ue/w8RQKe3XBttA3+kI8g63xXaDPQOMm8w
jFIVG2agBXDbqDpeToR1/FJEUm/KPQAJF38xyZd+fu86vGsdWyp0rurpj+OjDlhA9l+tD2E1eocX
0pirhPhZWfiGORMcD5gCb7z9DRFOi2BaLmdkMKIOzNPnDKl38npPPTjXQfyNEXKbaKxyqsC5bZix
CvKCVo1xrzE8zvgs7W5sJ8VFJaO5+sLUjgqmpUfXm8PZKrx0yoAobE91qi+wvUxNRokFIdTOzxIH
dsd7AIENmeugfhx3uFNiWPgsL6mMNCNGcd/myKobNCRvYAb3WL1fbPqI9qEOfvBM/oedVUjzi3LV
cAI5RbytYsaYLThDX0J7wTMZ2YdmNqOMWjjURk3DLK/300+UDplRS6gRPike4bn6qJwNTo7W/7ls
dkBvsq5tXki0HUw9NhJ+Un1IBpgeQfbZwAzfXen+tRcGAUiHriYQuEbpu2RiItW45h+OqZmytujd
e7ErSnBpZLndLrcG2Ek9PJY/OVvMzkBaN/l37dLk6IVdJjceBBTQ8URyu070IAoa4SzlzUvwff0h
dRto9hvUOvHpmlM9QeT3ooeNT2mV6WPAMncyuWe2qxs31WAn03Qs0xLWB0/VCtms1g31RKb0jTF2
mrXg/ydZ+fLAG/s4auiXfozidzSEIg5KNYVi9gCjZBVAAZ+UcGMRqKGcqZnicVn12EjIF0gmcRth
0epMQJlz8hYo2H04S7aogjFv8ylN3wCLOx6OO8in7x0DWcyWEXcwGCwyBBLql7GSC+zUl6IrbE0r
xQSxVfSvLekhGcegQ2XYt6hb1CyC7gKYxFurRbgX78D4J4cZe4tahOHanSFSJ6HhwlyVTdfRQGNq
A8J3vfG8VAfqwY1o03NZv1YnLLXhkMoiPGh1fwN2u6xAXhsoaeTpmw9hGPEQRq5qKcnxx6b6wiPT
0Xn9mwrpgyfDioq8Eu9cF1vBM5gbmkmf3Feq40HPdutW+snql6d+pZuxYZ5c7XtCJD9xR29UShvh
J30JBdGpNgPhya7LSl7vy1CmbjNrQWsHqc4f/N0XESN2HDr3vtEOWU8C9WfuFUlhwInA+jAcjL2E
zXWS/xcF223JRrJWJQWAOJ70DcfShLmeUHn9wJ2ufl+ucHTGr6tERB5wIlMKELBRxU8/G7ZFGG3v
ElsnAf4LYEz2PRi81srmorV/aJrl5WazIyll2bmzCfnjQEnT0O0ez8wNKJIqEd09Y9oRvcgjfb1e
ypHWH6S5rfJOFxxwqeIEHO8dV0Y6897dL7yb07DVwnHCHilMAqDN5T1f4NS4JTL0rIuNogoqfIaN
SuAnvALz96LE3MH66RxjXhCxIIXP0kosHE27+hjkKzqEyCKbXn2rJecO4HcNNboy4RKq1BkabAAP
kA+PqC0s88TRZgNruJGrIwemzRNA9NI/Ag8X4G23IXpuGTiWz06o2HTDg3zBu3Dd3oLOWG3m23vK
rH8mXbn6CSRIaE7wycwVrf9AsoHgksK+RnVndVUJsYX2d4zAd84CktQgz6gBO4FS6a0gA6jaV0uQ
YknpOMM9xpXIDN2W6/B3t2rUOnVMZYcC5CzOAaBZVIO9oufubJT/iwY8UekAzXLJZGWmmSkK7tlE
4+yAVQz3Dhj+RxtFGiyjuAdpHvPTnqaiLi7PunW5pzuRrtAZnFvk0DF98vunDLh2yMdkgsxMCJlN
TMSIAYZAH7f/8aUBCXhhkKZx7gk6urF1x9+aXALRO3GZvHNe/IlY7xLdkDhRvJxRsdsqnPdlzQsX
ipVFNGjp3lg972LU8XreA5aytM8pamCV5nGo88iQMX969rnqJRCl9foiArkRUpAq0/3A9ERpK/yT
0MwIjdhQ8vD8PtdPID0uGpvmmLhklaOY3NXX5GA5vjD+dRcC2cQVoNrVknrYJIY83wua7Km7uM4t
vYY8US+CLzQ0Y7fopmWV0UMP3/13uoUg4HlsrNqzHRD+4t9B9ms+CvSx7boEJVZxRqZS4y4rxkYM
ntlirKD41oKesoMKBYHgZ69BVNPSMmx1JXKPyA89wvkeJLEA9BaLJCXBmCltNXvOUk6w0H1qf2QX
+0vJ6DcJXiqCQi8e+PG7X1YvfAhpAd1SY/5iJaQe1oYcO7PM953n4X/3XiyjqFYEVJvmThpnAe/d
l5zTnn8ayOvXOLYJlfq4SdSKEBQk/w3+DijG1KC7SHpftiXGAkjUbgQkCuXFgQuKuU0i3WbolxOl
OMAsMQc06CKsJECJGXh1qPXJZgGGNeM60IZ1xLgJXZhDla7mDK9GmP9PvqvwRVlS8BRTRu3xRYrh
n3D3SunvIUtFGOR9GmJC9y/Sd0/w06orEB7WtwQvO43gUWEpGnt8mSegBym28mQbv6cJbgECXl57
EzrHqP5yRTSKrf+FqH3Aolsyti9Mf0Tt6ByESt8nlF6mAkvgx4BO6L8SqHJl+wSszbJSVm8bA54l
VAoK0PSUmaj1MyJISU1+oVIreFS/fIP4kyI1Gua1iKsBRRfPENvzGclwk/q+hNp8OzTVvYwMOuKr
TDilpWV2e0r5ggJiA190tpEqiMtwRFOELTkuaq1trbTiybqw3ZdtRFSbaqjzyHl93W96ACE+ITLy
eX120BItoAK6pv/dvvE621YYhl85/qCSj8hIWxVPpINn+vLtQwq+mBne9mDbUum5G7HDTY/RCyq8
BixAkOngTH7VSkfh5D6HCJ+hm6o0lYBOEtcaBtxtk9tbAN7WcvKvgOoymMQEgq3LhXGZwMtkNDDc
VYGzFBJtRajzZtAWGzch5N1sFzYD8PodiI4jb8JajnhA9Qjbn5uCsqIftHFH5z0Ef2IPX5xdSwHW
LlQ3IxNFedvJUddbU5Pi8fYsNzZ2d0oFrWSH4OhibauMx83xbv4YJqHZZIHubmHdwpnNFWVIFxe3
3gxQG0N8C2lrU8fqFpgXNa40N9xXHZdrhleX+rtmJRj9cduFNYxbgqGKNO6ycbfAYcz9kbHOj2UV
UTvsBjXhXg2j7xcK07QwV2KZNpKHF8UOEx1vSH+pe8vvs6WVBueOJm1wTEY5+Oro5yGF/gmC7iqJ
rCLZJfQTJvY3b/uPBePZ5O5KPM9R9zqojvwiJKX91YIcyMABAhWlwtdQjhYxSSbciu8ILW3grax8
6RwA9E9zmWqsiVw/0R0/x+0oHEvJALivckdLzTKMXpYZp9e3Rmg1CBdY+3CjUmuETBjhzWhNiWPG
/nmcTFR7o5OnmzilBMJyfyYeHnrfDfPDNX9jCYyg4gXKb1EQqpKUJo+u/A4rYHML9PBdW/DPOgDq
47nRLCVmbBG4vonhKIWbMofXAJN/4C4hDX1VrsFFXdqONyDTv/BYB5iI7bOFrhdPIvff9uWSNjM5
W5glqKeOeOu3PIqNo8OQe2iJ0t8UWyWEvLlQMxO+lW4ZZJ9pbAugAs9fpoQfJ3JDaTgsywA9txCB
Nd4TQ6BsfbZXxz9g5gWIjFQMQJJsnnDQg1IyyELx0eDQiZXrz8O8tNa0eKAy07wQZkzipYcTneT+
azTV/OquTOuTSLbyY5i4UHAOGtARQwVYWI0jBnjzfwmJZeWA9Gi9F63+mv9g0K1/ZDwcwIa/RBtK
XpIpNiynrxI/4lWCSPxVzTXzlKck3lau+6yLDd4IYAQFsdhZM+zUiZXE1QS6EzB3+ZoZs1MIHglN
tLhRZwKrJCjG9kZWSqkgHcCJMPTvlppPpl0FVyy/jHQc7wpld11708lbjVAcqv8u2cvOwHJ4iVzw
D6HOzr+Ud5TxgmzCzW17/o6+H82Xx4rYt630TilYuEK9y6B6F6Jp+QMTi7u/WP65q2LSnbRq1wCq
RxQngUcXUuX1g6VpKTpmnES3/v1rJlv3Hm9EBa1hnU6IjeFJGbxwrGSIVOnVr+rRtEjuwGZs9LKt
0M5I/J/2JrrWgJNHuqi6YV6p26bcZ0AXR0hjp2W3uGtvfgXCki/HYORVd81wdd7Vy07RVu00U8tg
WBX1DHfaB2PGO2m6VAFKzjBoev7lf72Q19Qj4DmFGPSFm6Fr/uTbGuiPOqziJeegAmBbbTWuFOsz
Jnmj9RJADeLlHf+WmvepU3qCEZnTRsthIhoj9CkOCKsdPqnFkPzFtWskpiNncLva+uZNX33A3QS6
lCOpwLwsHuM0JoljLei+RsoBSdiPDebwnBGfErMJT7L4nuKUbwLirliKQwPOa+Y+c1dkbviX94vj
G0V0iaS0VSrcSevebg/PQtV5gPEcwsxgcbI5nQYVvPaQO44n/xTcNSJbUQo8i6VX8TfSisF3WLKp
FNQu0R6+VdfTWQaxk0kB0aowyHsnLdvfqG5L0gSZSJqjj/CsCPYFgaagTtNz+y4UYrSQm6cRL57+
kY7l3eapnf4F0yKYd+ST7AZ+6DEc0ZXr+A5hrWCn2ft1gfEN7jX3iyribm0VfSvQwdjY6MDmgnKQ
DMOX4hzY6egdHWHY9GPGz8LwB6tkJwLduA/M3MeiJ3fa0dsLfENSJKFAyoFPorU47dvct9rIC6Cj
f0pKsWHkOLRfrbhAgYigruvgWsnIfYCan1qVGAFpJzA72hp7AAsMBrpcWKenKzBMeavkGHi0MjIR
k5Sr7s0UW7/0OInh7MQbP9STLvHsszv/2dEa4N2NR4cc1bgqoGSRVWjd5/ZLThOk5YYaVvEyHJ5D
+ErDUZxtHsxWQDGyeNbvqwgSFnbJ5tctE0+FBf1v3Eave1Dg1LmskSjslDGr9j2s0QPQn+lvhkoo
qAzvgDsk1gM30hg38wa4RwIMyajL9mo4vsfAXDyxL8KexzKkdBGIXN2aQqrlhIjbIiSW3Mf9X7Ut
YntpR8UuVPBD+mL0kM/uioEB5SmzMJ8/k6Z4WpFq6vc/3swzTcOv1SI702WWwQHHFAKsi7Zn8K8s
7tGIHIBCV6aAUaZ3agIx+nbNa9WD8v+p83suKiuPla1flx6jtlk1HbRC10aH+zLJWOkKV1kL2CsI
3hErZtgEt/tFgCw3XfIG0t20IYz5Neio+wnOdPBOVq5S3BCw7P+E8gJmz+J5+IFOhGZgGyGFmvxq
BFy2U7I1zVrc0tpfflbNo2qkRjR/jEPQX8CudYevCWl7QO+tp6M/QNS0vRErhTPwIlnp2bkcjeSs
dv4yz5aNHlMgvE30S0C8aY8fV2Ww8u3rZ00XRs5gD5SYV10rAdxiGgMFuZ6+WrkMnypMvEk1AOum
EVMCWrKs/KncLwVpL0VTNvtESVtkCoibXOZ/Y4AqilQtjgw0+riMypZ/M2hZkFmVStHMwqprFPpT
sR18KfhdpLWKAPj1U+DxygdE5Q+n9op6vq+E25s+V/3oMoUbtKSt/M7U2S35qVUcBK0Mjiun+LAp
VJTCkhTdc9WBRFmsZV6zIXpsvLqgobpyw9SFIZ+Wy8IJQBfRdx8L9nIegM/PH6kVmG0izE6X+aYt
My9wqY+4anbsqSrrzXl/WW4zC/jsE0hVzLJjf/LibEbVjLPPK9CxCsYI7MbjIzl1Ns/ifULeVxM6
27CC8/xdAC0JDoFeSUxHwo5bc5j0TNj0brE4QRGcy0yyITXlfhFVMlGaAuqQwossnNoGcBhJtIZu
VChNY6eEFFru7kwAr2KI/d/+R95h4/tKmnpNdI2taaTSYiUvdENSpaP+LW9wrKS/ktg7fXGsojo7
psmFVdTYvYdBIpZLDeQvIaRDPia88bAICEvR4BIfmJEKCxtLFUN0ShOrlWz5Nd7wkpMIVLUpWAAL
l03PDnHlV2pnwdMtQ82X/EaCnFHseAlAakr05nwVC2d4MyXC8mPGbDrdupvtnphx6uJcHIzy4OBg
ESrEsN0HDn3z77AlwoaiRUUpre1s07OSixa6Vesd0bXKyee2FVz6BnGFV4zvc1o3D4tG+DlR4SQU
Q8oqYjz8bwuqNVoGtxcPxX5nZr/66P9E/XGTZ2Nnow+m1LZqKI8hD2lf491WuwbU0ng+8NQegBrP
NaeEK60VZL57VVVraWXnRLvZPOqGJkxYmA/c97xhVHMiHKPmlutP8/8qu/DUC7mHatx4gyBVOMcj
02662udhFUh1ujE4LBgkAyTU8/aUsu7r6z/Zs0cY2SXlSg2lKxeFNIkKPgKKLL0dZnyWw74To1jS
9MzCA8QeYDVacacojHQRnW/OLMptb3rSTNmipL6rlAQgOPwwRQwL9yETbYw13J3rrM0nUapdDXxY
tyhtxhWFSWNWR96KRJ//jWqNLLV+XnyX45fB6Z8JaUj3FyuCxNV9rrhMLRaotjMwqAPeufRp7lyO
OR+40eJb9xFo0+7jTHl0JkQOndlN3WDxfQ0VNJradtMLFVGKIS9xqnnFK8mcecbJ78RAVQKF4X8N
a35lScVAknXDJ6dZBJYd4HxiebSGeMcuyGItlnL0aNMgA649RNidmn2KYJALlI6fz0oRr96LV+ms
dbljKV2k2ayNigk+ZyPOthNU0MWWxKww0D36ycdJEh0y6WSbDc/laLWjbHU0bY5sa1zR+qipgzvl
U+k6sdztruqfTT+GWIs90TklFfOx0IWo22LYkcLF97aVKY/kjg5NfQhtVkSisTIWk6WbrmXa1BFR
2XJyB8yUth0POqNztyVFDnJFQVQWaKa71sKYCwG81rrDxvqmAs3yi/o+JfKy1AOAHHoJD5VizNNh
SI/u1j3GlC/HIjM9Sgkn1N/O2U02OAn+X8HhPcGyh2xrc+KtYrNBgVCnTa/yZTOX7/xctQhhvWAq
caxXwYfoI9RguiORl3Pu1eltPq2v0KMwWDvu15vhbm/C1jFsmRGNwaLpJwv8ZoCNu3bQV3Y3MbjI
9cAcRGLIhsTn4mbNpBlrQYB/4f1xMPtVaomrJ9fBpe9yl+t1Vg/NUgUFHrWzda4TPU3liSG4CV3h
hEoPWGToMQ8WmQjvGP1HDQSCZrwb9isG5fY0Gwg60z9p+0BxUZfVSWOl97KBu54YTcYHperL+nhv
1rj4AwSgD1ejn3Gh3yZLi3gpxIYi9LI4/Y5DXiVPT1hbLjYYZBtjbBoLCBYcXY6db7aV4cYfCdq+
LfCQmBHWrcpDMe5vDBLGQ52NiW27pdbqM8loWKShwG17phUR8l/yAOaCQo38K1WdeNeedSGxZ9mS
UkoK9ahf7BHncdh0nNFGTOkrN1VWjgOOP0QVATpgHvnHG133iDlFj/hkvG/AAnE8nN7UKQB8zSSp
wo0sOwXWdfzwKDimD/2zt73FbtpX4wcKXovG16Cl1pfXM6ZHHNWR/atbSpJmnbO0d9YJTduR0PSi
qbsBuqAeoFTCMDBXA6FnQO0ZMM3Q495JeCeN9VYSTsocb1+xPw6bsb1O76TOyNFV6rrAYTNJzPkw
LhflQmXHd2ll+CYJRe3jh9d45Ife94fajSM6RTGwhfw0UPg5PBCP/zx2UXXCNvXUhSeYDiEfj2ca
ekGab92atjs2MbL0NIN8vtSJf3g2j/TOFf6xJCK1GnNUHCd4CJ8u7ha0NQhHFInVZmgpEwZEtgLM
Fyzb07u1ePIzvIklcWYaO/2V7lWYUYAp40Mdpl5dUzsUBI87F8plAQJ2N79lCqqLnOGWsx/mLvIH
QBRMtdh/fhiYkQttQ6smyuDL+B5DG6mQqw+1U7G3pS7gO4EiqCpSfn2hXqDXVwhsHNqi3lalBiaI
OMbCZLe4+CA7lUO7mmaZMWwkMnn3ypUhNS8zTNMIaA52lQlSeX49UsJaa+ipPoMtwdgC5x4lP89/
VU6+rbc9mx8Uzcf3cHPpS6wDCviVE4H6jWOqzLFIBuJ88oEsghvL+Py2m2uj4ty8hVfYNGnkKZcM
lbtxR/KyJ0tvk3w9E/8puhQkC5/QAfE+xuVw79dpKR3WyjSO/QXoTCsAXDvWvZW15q+DzlkjwQxc
sMJK4G2qw/naRZ20kk9SYnN3Uj7Pf4++U3OGAnrzGRKr67JIU3qKAYbpKfvVuSFqJkKV6YJDPCaD
Tql5bhL/uRiv1W4WEAUeUjVpuG25VRLW0zr/NGTNE7+RBHhfpfTBbAgxtxD9IsMo9U7MdCMjNfVU
x5qpCBfLPoyedxXmmVEbTGDebnCQ1OaMCXLCWGE6GpxIAgM6BlHwiqf7NYqs1PWWomWcH9obOK1s
je/8Nnsvmyww2ckh1eSjXnnERY8m8O/UsUBZvbumfZ/Q1Cj/TApVQecClm3558ECffXDk4SHfoeJ
GKfC8/hzfpC+WYI3CcgN/9gGmOIS97o7j1fE+Eg6COs2HZxA5WeIWJexQBTvawNSFD3gOy8OzVoq
aIN7vP7D+MRLLO4Hum3Xtq+7X3RPPd0jPsuzcu6AcMwIkIsOzsa5qwhkVcuoRwxavGrZHuRBOKnB
C/ADbsPmH1VOyNdbImZCujMy5WJptG4gU8xgKRfC3SwawnNBH60EVvdvis3b+ecwIXsKDxN2/cXw
BGz3YoyzK1qwj9dDBcaK2wxoVcdthIuMkpbIiMDTiIOTcjLNoMf625J2QAa9nYwLySyqZJ65u71+
Rh4vnIDQANl5S0NffMVnrFn25xIn8ph2Kl0u72tsyNSFh8gl22E2qbr4e15iVGZ+vhWykNJqf0NW
y2t6RTFeEVID4hxGOIV3mTMdXccW7uuVChqfZLioY+QEf0unL8KVFacF/kx+6xE1iLHdJQXTXZr0
EgJh+f9B28TyW4YwQJ1LetCcqt0kNiztrp0FTpjLw9+gMFno2eodvnfmq5Tjaaetaw7xHEIWAhhx
ILjmLBdW07PLtFk3VhHbuUE7QZrNWABKB2LNCmLvBmJzEn+XpRekdUIkTXAdnie9VyjqfcCvX4Aq
622I5lN2eNpxOoxCGiYTwQIC4/VjYz7MhwLOdNrjQdE1EPZW6T+v6oM8F2hN54bJ2Mqcy+YOE0fW
bpu0WYWjvJOesPH5ndjrVHnJSTZVMddETgr9xctkI62ckP7Wijq1LLoi1AGnF3csuBd5Lj1El72q
U+oA0pv24MOs3CF/1WjAdHRoyL9cd8wYP3xaZlwgEm8J0RAEgVtdGSy5/7knshB4pT+GddWdlibh
nKMV8QXwsT2kWh2RLhj9msvDRJqwWasLoYrDn2+OCY7IqH0lAi8xJ/2iI3jzbWGlNtjYgYDnzrPc
Jl1Ufs8BaKWMGkap8eRkenPvFuJRG8DYW4veU3bjvnmmFDe52dycqyrK+PIGZc0BbC4kS148ZXlF
x2MjpEp+W2RGsBDVSnOu0iagVoWYaQKz9lj4qFKqxw8Y/gUKxexOs0hTgmmUjxiz+5ChnOYA9Ute
vHso0hhrkWctGWe4hh5otH9OxgYeSTWTJkwSWTuiyaluMNi88xED+Li8jPToprRPgw3l8CPtmwgT
EqsNFlH2RATKXjub1xmHqg5oup9UHQI3NE28SMfr7wJJ37D7J677biIA5p0LFVap15JTKXSxwCrR
wDTkGpuWtZHvvwKv5w1g/6NDtfxD4WOx9Z+0+TC5Y/EZGmxGQPFKCoEpSj0dsm+Gwa7cGpn1fZr0
U6S7UduHzoY+h/120UE1xVR4nB/eXEQgJcG7L3jE7ofk6cVrEPZSsVgTerePO2zTQEHydH5T9cpD
UPPlDIU7zx3iqkazb62ZnLWyBH/4HimqPQeVCvwaqTnHTHI0M9QU27gQtlR2nLhfJbOmbr7r6tl1
0Dx4YCl3GverijGUDpAIQCtyAslDrAcR+Pt7mIZMgTrNpfAwiRdKqGwzq7pgZKdwOWlvyEpthg83
CafxFj+Xs022EBBr7r78nBBTWUf5Q8GAgaDOn20mF5hNnMuRCs9aqBV0Ra7ScJ7zFwS2ap2j8AXd
dCyEvRm+wQ2g2h7d54E/Zza22OGwoYWVfmfcCdItJrnDfYCwoBH9kHiBmVbOfwzoOeNMZZ104SNh
9S/S6UZj5c0lvF6cOonEic7Nlht7ijBwL28tuTheGx9K+ZPJk/bFbzErfhKR/QP3XAmpGs6OyFIh
lum5hhKEVEQ1AceMTiTuWsuucApF/RkOhO16nrqkYRpZUMq6rm5pMiimr83m/THg+3CF/Swnco5H
5BT4qhoxKxB4wq0DSvSCLi9LA8nVQNB8YRihDhQMzkCe/sOaktXrqaCOBEUKSD4k3ADTPvgh+u6e
cv5fBryTsqKr1IR+5Q27l4IKQltO5P2EGXRyPZ1jJ7hOKwp6/5THQfyaFCc15B/tBFi3ZoT0FgKj
Oh1KBAXXSN57yOQyUXEjajOa3ZRRJB7T4/ogvC6d9Rqy1gP2c+NL9FEk1mMQBKVUl0PHZj7+TSnf
OfAJPA8lSRAT4fszoDisvmxJ4tiidDpK/rAd6vlpE8rg/57UwBtdjMYcS2rC1AyZz1qEACdxdoVW
cLSsIIS4UaNf3OnQGEpuPtQ3r0YfF+dRjaBIX6iYSwL54TdNwby7UCngQhbALtdAXwSD3+Q2EdmY
rtBt8frNgjxwxYGbD7DL3qRgaQCX3QOF/e8GZlXVCUe8AK2QzmXKpb0IuhL50S33/JlVhzQqn8YH
JKBYtnFtPm/WKWjHdqFZkwBF0TcwYb2JNFbtIfZl+XHj3EgurDsIThTY13rn4vaDEy6tQ21CxW6U
TYSl2SazMM7+THWMJMQWPHvKGTvKi4+EzLZuAiRXfoV8LFz19AcI7AyaUMQri0FUBkTk6ZrX6NtH
DtNIGipLPI2u+3DvO/1cIz3VpvrAoXBujMWpnBAW9C79957AuF9v6hl9Rt0qRA0KgU7uVMJI4SgM
EZHunUm1rvGo2rDCF1xR/nhePcv54a7T/O/AMy2W9ck7DebD8Ea0xM+CHPaJP1ym5mMOnQKUopYN
fmDQ8fztPRm+z94CUQaA43iTPf3aV/3RI9fEBr0+yYwIkLt0PqaIo840Ui9GkWnfUCaZ0+/X67gV
SazePSfZuL1Mwu6dPoo3RX81u5ED9raKlT8SmivrtwyvSzuUZB5j9zZjanQroSwZrWmmtYOFAM4j
WqJIkHsRVM6XQbDeGNvmFL5dsxt3jzdhMIIklqGCl1BSRAQmecvh0OYPJCzJ+GejAdwy7zeB/DvM
Q5pwRLeQ0gDyJaGMrAjtQ4ajbxJAanpgmgdbwwMiILYvxW2i7ZO6Yxm4QSUsxHTdi23F/8xV/rB4
xh7oBOaOaM3v+hDMaPHCxFyY2db95yVAeoXSaWFZagry1TmiaaWDyZWbNnoj6kr77OoehM1ELwJ2
6uVb9Y4CBVUGqTUq2OnjpTw9hVltCVkESjt5F9DcN01Lot5NZ71gD9IrNqEv+5Lz4I4kquSV9+jC
5v1d0wzRlyk6QOczbEnyiQLPpDntq+EFFzF9AxsfWcTbbTB1tvLpW075JJ5UlBDPb64PpO0uHVLL
AflP0jUvIi7sHp42m6YZvG8C8JSW/rYsvDttMBPRQTLuz4VOwfMmQKWV3MqfmU99xXMmQ1hh6RLF
4jsWhwwRHIvv4GTZWd68JuaAvRt3WczMuPI9IdBDGKi2aSAhrqKb3saYahPFHbK7ii5VzvyOEHZ3
98c67jGTfWNgZAN1BOykMrSzppsBREGnPWpdpoiJGXWFMFJT/g5hkuh96B2dU9LMg3i7X0/guBx2
XYZovH6lqqZmr3xHsRQ5mmlSpUujxD1gTEERXPxSpFi2iJ0lQiEto7qUQCMqRbBAomatA0TmXx4O
RHSZ4QUVDBdbvLDVK1uGz5niPhQUnbFp58d+pBIuDuxSUDvnMArdmR82R3DFCCAU34qjDxnf6g7n
LhJtP74gfzFWiOuvRNHOquz/wU3kymfngcL99W5+UJ6GnwPtJo/4S9+xZXK3FgDvhPhGskjnzldR
NwpnjfrEnX4hawzfnNIMg2AcPUe2inJCCAaAcv0uilJThIi1862DMThvu5a+X08ttwJrw2ay+SUI
NFvp1xeLWrliB96e7KW59fy3gaosl0M/CaQuERJ3sUSF3ec0yNn+aQo9tR4JPt9hrhf2RTwkxTVI
EXlHb0wz/zYGRXLEATRCPopdrLCslYyBLKy3UIIijmwEcKVnVZWpoA9YZ9HBcb18kf4Grj1Sbpe3
NaLxIh0IyxBOjw4hwqMZZ11iBAIlSIilQ5pQPTkRGRGukTtCI8NCFSrUOSqAIvCSZzlb1i2iHG8K
PbOb3ke5FzNaom0iENqCXmdalrBhN7oCzzVBNqKqpmynpWS3/tpuzDNST/kExcZQRXHoL4xHe24s
goK3NrRldljgyxiLlEhdjuOTGs79G0jWgm1m+3AB/KlG9LtCdg2u7C0uwsC/wD3T5FtDRouiMFIs
kExd6v5g7AmCyLoaQtAQ8uQzgegmIr5LH+6o174eyVXZ7EfKYZrv1WVwbom9GB1oiPF0f9XqrnTd
5YlreIvVdP9trhbgOrQv4eos3HmH2OqFw/0qj51IO5PBMgu9vY3i5D6EPQZEJevLlJCEyFXVtxvB
F3+TUi0FswoWcYaOvNfSf8ceCM7euYm2Xc159r0sO23CeCUd36UAlbau7Mx5HoIXhGFwz8EE6WZS
XEQRaKKuBJ/c5usidMmf/aPPpWCChhxDA0SpvfRWzIkvhD9TveJBv4kDTYGGHot8HN+SICqIDvem
GcapAbF0uxhj4X3w+l6VUHsKJp6cvTQu1hbI9PYOlAQy1XJEzo6LRhd7qBSHU5z8vkRcZRB18SMq
OPvOfwdh5PWnbSDNhcB3Py6rEO+IiT+Nv4cjxiRlFxf74R2Y5by3OiOpDpBKsnPP9QwZVdzL2OTq
Brxlj44APuN56GnUwPFHRh9sVUM+c6SYNuX5IRVbAzBtkYVhWG6drPf+0N/eD5nYLzLk9TXzPCFD
UC32f+lKn8n4WaQBKyJvayTgxxQmr6LVhhI6uTKYGzVGJctQwz4VgHyuN9RcO1uoeiCfuiB0qQGk
6O39/7CqEarg9ag3gR2f2KBjFR1iZetxe+iJNk7vQl/8fJSr16BfoxwgiGZ5/wbHhLQKJWqcT3DM
Pa1Bjs81KT1idKjnAfavQh4tHl6WeHsAz8UjCGaFT3B7Tyvy5KmQKksOv8ZRodOQOqbEAzXASE5B
tt6FS86xY62o51iCxpu0UK/CHej+NlBozm8S/zJz66iIV8cD4O2WgoJO6FW8WoITe6WtLZB6sSOK
76gyAI3jfcY92dFrPUZ5fMBfZ6LoC/YvJqQ3Rn0YmhmSxfYM+G4h/QV6jehsDx/jsH+pBdytu/52
Doudkx3UgszDeOvsNzwzlv9tOtrpbGUk400gXzh+5xBF37vrDBnrAdIhLOXvrxBlBZl361H6IFiJ
c8e/0zJ+pPrNYhv172Fap+56BQ9qlRfqvn+oH9O4kUsK2iFXm6u0+Lz2y0py6HcifjuCjje+uirR
kujCoucfMTu6wSOaat3XpqvYYx0iQhuYJ7y8340nD5a/ElFudTjgsaxtIFDRjFUSb9verRMjvZuN
cLzoB0mZ8aEBCKrzXvscraWQ9b+Of9ukE+vOfh3zNQFcyfth/vU6wTJ0oNFARqbkCM1iyLEYJPbY
qhVaQ8yE0mRFS1TwuX0RizUQrorU1O3p8i+gwq+2BvWSaSqVWdEF6W+ca9tcMmwvIxO56jbQtk52
CI53O258u/iq+SZYvHCKlInMcmZsYIOeoK32u0LVZaFsOyjatpdIu1XEPnjmxjKEMNKq0eaBG9uO
+U6pIvCGxt2on9XsdIHW4oPPlyarPam7hQXCNIFn+VhWrQGwKVGIbKN0dczlcexABl1tHQeZiohd
A+fA3m2YrydOv9L7VEvHaVYaCbBt5WJuWhjFOWgCqJIOlGjQ2REe9WWK+Mfu865FAtaVFrzeAH5C
R9/0x0rH9fulxPflsihRscPGiqtujTMu4xzGuoESR95Y2SJp0Eo65JZC8ajE1XCGDndH+xU/N1KO
u+VXvuvb4n/DJYEY0Vj1GNuB5PubtS+sg54BKaCPlgAGqXUM2QggRbH+rt/5XbK+Mv3NWxS26Ee5
LY9Jt10itV5XxnJ5L4WrrvK4xvINkLpLHm+lz2VrUvWTYlRdZWNllQPBol+L3IhwiANFKf0J5Mlv
NhOxFEWJIaBM6WmsXlpekxxBsrtN51ogVqhDkvrUV+qZ6ETJgXJVvnmFYbsVRJcCbxv/d3wUYfCu
skYkeQYF8sl/S+W2M0zYvjwJSbv3yBbhLbJqi93euJYeKds6p6nKPdNhB3WVEYaXMeBBH9HxCS1A
wLODLxBuGFIuyxK2Pex+MurfcPLCQ5r5jOOpm3dR6oIllj6Pd7w1qzeqDzkpxd2OCCJwpU4GaHT7
hMYs+nSh5x9CcKON3SJzto9dW3LnsATMvq6wFJvs9IUfsNfGAGIDWEHk9RKj+H4KllLfY0+mVnnM
AJP/3AF3F7spMe6SJ9x0H1qB+MU1UqfJy05lhHRkoPkh5u6ZWN5s8myZUAOqnUGEN7bfFCtMn3xI
73o6BjqYdFuwWo2pzcuaLEg2yavIVoXTnw8EgED0LYecluQrtbAmtTgn6mgGDLh2BUVoGMRtDtx4
e0T4S/Lsmc3SX/8s7FvwiHXC+YFNTQwnx32JhpM5U8ITheT1GjmJzsliYNU6isAzuDbWucSIoQ2b
4iEjFKLPgjUuHjc/GxZHPoaOrNDCLehcKL49kW/wPWqpn8kBEC69QfyWvItVqrgzVesh4zRl6Mra
PNGdQ9Pvnn0/WkTFGW5z8cE4ZKet7LdqlvezSjTD1b9hBlDsDkzZmAGpLICOdHHZMlinthp8XjoR
WNdDSAIwutMOa29orHC/DtQz+PVGKhivDblfpF82SPSOxsJBL/oaCJ/KrptM/OE/S6AHp0jUCpXh
SBUjtYFVNdM5oXL0M9jEE4/kZx0SdtFMLi1aoulJuhuJdNckuZt3OZ9ZsMTZkxB58Lg/oAUJ4mYF
O+A4s9aIselTjQji/3kblzvkX+IKi9YK6/M/Hbmst1+53XoLplJt5fASFTpC8yaCTppxa/U0zbkx
31sFzAkC/YZ4qJeqYMrbv5fEOEaA3gqwDomDUjAEARgzEdus3JBAvpn829edtqgg8T78OpvexLiQ
qDwEV0RJdVuu7jp4w5OAAK1UMDzXQk5f5fckzqz0KzJwZ2YKJxve1IViCK2/srTK8/MmOYbgPjIk
n7+B2BgZL6HRzS1wo85dJhHNcR4D3RFSeMKPzcjuxyHBJe4TXyemcM4GfC1Y9XSzrQwDzM0BNSQG
RBvQVekx07h/eJzGttMDXtMwc9BuTUjX5TEvV0ys5IWsjqyZ+zn6qHggeCWzRRxzdIqUO5WHVuRy
+Xh3cVuKPcvjxkDQOJzL8FN4b0dWSMQp1GpTscmYwjX6kpeXSgI689ioCz5IMJrQmCbYJrHJou8D
Ej6PrdXfK74WunrYhy29IQ1+L1rSh2JxoTg0GdD6FdWCYB8ildXcRRwarHjpttg5gCUuTu9mlm+A
s3/qaAAJiLE9Zesg6MLIaDaY40R4dYYF2+XzEW0kFKdF2xgM7sZv5OOgqZ4kE1Yz9R2NiLbt+8ZY
TrwFP5usPBBn6VBcOAS6nOOXc4dtV/350e4Dd9BcK7OxVb0OkYBKqj//ctXxJd52+A0wF2h5BwOp
ThqV8ea8Vw3CNj05XYahDx1s6/8P2ytLkEq6Y2E3bqJlamXix104y4JBC8v81BEqlIGZWxt3+ZGS
mYg+xLe+hk0tGoBYhpXKTy5qWdOyqgfvYh5OGilj8j5VXfLeKWD/640rr/myCLEDsLsKkn7wYPBo
O0sqFcKs/JBlbigDybIfk2yqCp/h1yTusiZ0LK0WaB4ZToDKc3KUVn/P64NQK5/8wspzK384QkvY
yeXhtHyCn+epUMTjsPijtsmq6sUzfw1rP6LvtovWlrQ8M868cM87KPDTS6f4LMRfM4LKw5fLWFlg
AHw15mUxlKZrz6eAXycjuaQoe3T2Rnkg2yRPgzy3cVXcdIfAEYFuV2hd4Cr717gItZ7D9OhhscJr
yuS630XJD785QNAXYbkma5Sn0bG34o/bemA4kSw9sxHSExjoiO0GJwPSorTpstr0kdUAfjok8BY8
3N94xzBLZFy30ndiRV0zeuZYh8C8B4lg9r5TAzn1xQbIU3eJTzR191JgV0OJPVSvt574s0BlciIz
2nDffLFR4cF6cVYAnETmAE+T+d4fvAGqg426LugJ9lkIaFo+LK33nwyyW9IUj9DARcQQ8MBNpEwe
nZxmQng9EsQqyEA07FirjXGcKKjA0OLywj5wSU15mXf3DN8bOOcB/pMEwcLacyU5tg6vufvvUNKN
QWhO+PAJ1CRffyFIhzsJj8QzQpizfvucBccWGppN+fagtWpBCXAkHkYBEln38yqrGAcMdxvn4pR2
6mdWGl7fDuFom5hQxU5GVi/9FbeEM/Pj/b1uv2eqUD+YRAkVvn8BUr8Jc9XPPCk+fI+Eens7OMVU
JgKp9AFbyxZotyzr75QWb1FsKQNhdBxYvTwVb8pwjrxDkZmKntPXSA+31+Zhwy4JrwNRNYCfM53b
GierDJU2+ZGlr6x3oCggS3lrUGPvi3v2YVSxVe3Xod/cL3FcPj5tT8vIsfHsgrbx5xt08BwwimnZ
yLtVsNNfyUwMS77KuW+dHfJlYofZpZacDdGrum7W3ekdRwWllOXOhGlxC/44plWpzKyHT1SiC0/F
nDPaDrmYIH4LAz4vV1OsTq99fstgvTp8oBtggk1HfKd7lMgXaB8Qu/mcdWUswuVr86tl2ILdGl/t
YcmIXrQVLDbP4G8ghFmhB6s5YWlKySKqt1oA7sQSjcV8Kda19hbc7phl+pYVDegjQ4CP2tXUe0fP
cLU3FQr4eQcMG3zYjtmC2mcvFqglX2Tl1zPwRD6FMGbHuDgZH7ri76Gm2k0i1AgkTwTXjLQ9MK+N
Dtthu2KAfUvhtvh9E3ecIIARgT046Iw5AaKNrBuy6diPontennxNVXAzayI8dINuhyKT+WbSxiW/
p/IRiY9G6aB66UjVUSnSpGv6bYvXMHoLQnOR42nE3Ktc45mm67MmDgFb9ORUmq9n5I6p/ZVHETjw
S7dWZgYHC9PS3ORXv7ki+oWXOc9TFqtpII2O03gYVvIJHvQ/3qqBQDKohi1YMgjMbw31RQs+GF/v
nuWgw2g3Z9NZ/TAn83cNsR3JaMrL90TbB7mrIV125kIwNWC5rqwDPeQUaCpe/6nL3ONpOlqs3ASy
NPcAKfbKnRQKVLZVL4I8BxgnLvFFwduqsRfb8MTdlyEkaQodjvI+/aank1l58LG+7cwOXMVIz3tC
wP7qn3+fXyMMNApdkYjgkPYoQwbJ0OFfksGPnMGIZCXul62mwv0SkiMs/ZdNKZg8hF8Le+u8J186
HtcFA+/8XtxeabtSKt6GL4xnbMH2v12JtHvVLFsRMqh2neoLd1XJvu4mwDo3YNNkxHksV87LWNZX
pIKn7fbHldQkPBH0GLNR9UaBL59k75QUSZ2U0neNNwQAi+qpYxkjC63t+OPnSRPj7KOam9KNKvIO
ivmyiEyjvgsamLzI4HK0eMrGpQ80CZAeOMLctnGf9TEI+2GiCQr9y+WzRGGDZY2gN2FMYB5zd9ue
9iXIynXNuTtTXgQCND6K8ysccEqF4ukjbDK3sbP+7HAjqscPd4U8MikNaIYWcxrq7Obn89eM9rG/
IfBxFVn8WwlUS17sljR9zBhjDAH7VOgMjnZRDCXYrNucyawVgPl0t/MMTDJ+hyaZ6VHfRTx61Sda
jAxcvKpT3c8MzxF+fek4UjYfBxMxPpcPcoLtcB5RFsIUhDrBaR88NjuSFBtIQ/Hd8+YUV2tFpCoc
7gt6LUlRYnOYR2hW2VrI6KzJuBKyLNMAuI7JzF3skWxoZuRdv2yMZkxWgkF28amPxElTm6xoQnZy
a2WNila+OQwe93dGAJ717cO3I4q9VX+8zQQngOrhv8mq4/9iar+zxic23iyb79YEY1kMZkTiJb1/
4iUVnEZuPI8il1BRf+caIkrs4W2IXjWhgjGihpLWYjsLDzEOp2HIcRKY/K/cMqXQgKvUtgIVF+cv
LlLh/1oLPSinZF8iGqh17h3D0v3QbNLOZp28MDjM6CCitk6aJlHuxAz6G5byj4aqBvG1M5CxDgNW
99cZmAWgizWQWpchXpBTWENEfEY5+aNxX2RMUOrDunQND1b42pSW1e2qgnniI1GOiOLQeRftfERx
3/4N00GIZOAx7e8gM8QKNTBqXXyWNHvtWd4am4ih7kwWXaf39jdAIHJ4tcBNq6Qo4uqFtSQT6IcH
e9q0RWICpFswTLXRnZ+nUsPSbDpH4PtzZYnKVIxcZC167w8VSQiDu06QBmNx5M0J/JVT2K7PZC9o
FZ1mDoWt8RWDsujxEdsxHK4klSaBgvBQZE6utfRifOdDsmDSQoFvBsT3/Plre0kJA47RNHYsMzav
qeMyUSzOh3GZtQrSs/2O1X5+NE7xDdFi2isHn0HDfmqgYJ24WdYxHBPhrO/+asCYV7+nzgmnuQ8c
JqVyTgJyMg6xeyeHgP8SWrx7RtHoDItiwJ2Od2Gi1Or/6sDPfOoihj/ba26HAE6BnvzJQ3YwLIz9
HcF93b6RCPzjXrDeUywtzGgquul/0KmjOs892w23dmishSxbvSUyRE+WSTbc08ZtpbQCyrGPa6Z1
rW/O43idtWoHH3Gi06O5s7QiNzwKSi9RA4aaTG4Fj0equmdwBX/MdZ3r66AS1UWRXVv1IRMSkbt6
QCHqBV+dr0cgqBjI9gdhse1QfrCf5X+icw/UFnyUb5NDDDtybiNpDZ26y3OCr/PSRBgchiYRbeTg
kTa3OibEDQnb9RMfOs4IitKdcWjrSbpNXjqx8wLIs4Wq/PW3K93k/IEwB01tDqmH00h6/PW5UBRC
pZFYT+qkNK91OQy8Pt6VnFLLhV09R2XmFYo1axTwUS1tL/i+L/y+JBqNodqXs4eLQLfhEGnp5a3k
hhhH0Dv3ej7r6gWb26QV8iG19OvZzeWRd962DE+zMSDT9fO3K4uPcgQrMBb5PMm94an2a5feDjHh
VHseC6yN8CMVBXcLfjIfme6o4URaVcC6LVnccUfaYrsFMDMWHL5g2cEnen69N7gv5F15vMM2Hae0
No8YBRDQj8GHBlFZ+nWnLES7YlmABukuUDRhGr5nT31s6lign5HD5+IACGGamjUrdFIJ8MS90POJ
bhWx8Cog3081AQYEytDHATyvvEguktNc/Um1RMd/Uq869JEHCa62fzzdSkGuwSStBR9fr89hPoQn
ol+dwJPHE6azonpM0P83DxrYksn08tfHBDC3II1var+wsRrd/iR4LbQcZlPAYVG4tmNmGx7kYuAf
q79C/ul5OxIuIru5JCOMxP3oMQ1EWvXSTU/cuY+Po/kFyrAHsSfNvZ7bExZHmF+h/FqWT8wZ2IBI
AYmS92u6A/T+i3Lzmz/AdYDYKrSgomr6bkfqkJOgsL5RHZziIhUhozd66zkT8yIUGnf78/PpvE1e
sF9JJg73MIiEm+y5g6TxgI5RNsOKz36JhcQ+HDVFcUtRSheV6dADOnJfj+88t93+sIHGJYKd7np6
cUKYVNc1n0gQScVVOT8Y8gjlRb7n8kIsCSbN8OynmELkf2Me4zMjVRw/X+ZkMh4fK64XqWqfKw77
58OHZ+SXlu8zghwtELPnwWNZan3YXS79MAPg9iiyWvjaBJc+cKzlLu+svj5fSDxTuXDv+M3TzGlQ
cXmLU9k6HDGef76zCmdsoUhg/43PcQJQXnAArlMcmv5BVPz5E4U0DPSKFkMcTSYu8dTMGEgn4ukH
5YFUH9BgqPrHgiDOAjHPR0U6XH9Kxx7On/b/fW/O4kEL75iXCglRe7uSRyvWi2NPC/BkJAvgHOWy
HJRMohViI4YOjpN3hZR3SMDpaFsVvRr45rA5fJ02TVoRag7pzF2vWntktZ96bcJnxEE3DLlq9uI4
SGWJzV3hqSArVqRpSpr0J+Qpls/zBDZ4myytErufBXgXXc4JFlLFOSV1h//+aySzVnCNrEi4TzKt
aJQ6LAnfy4icJYBDKg4LWYVh+YSr/T4NpreKjRs84LtQvQ5rTgM8io4BzmlwnBx4ZBAGml6AU1hO
yXQs+1HVZHImhe7pR4P+a/bjJH4sL4iJgUf5GHaS0Hm/e1hgYcInFLchJXZgqNgKO6FYtgTlj4RB
y95jNd4vD0uYlpvx0vn2sMFyfZAjw7XFLiELYmelSISbU+touQ+XwQhcfal7WXIPphZPDEN1d7i1
qI7ulkbDxCer6Rcpg5o0uw86DNm37VmHetwRjLF2gUhYfBmD6CLn+rZsvQRWx2qrsaX6V1ifZdYS
Bv1vRKnA+v5ExtWPilXReeBLvcjlcMRaAQGAIAV6Heyu0YBg7EWMetUw/83jcvHRnQX2QlSb0ZEi
oXhQHP+XGtPoNa/4UG5fZNYm5BH4cEdYKg0MHpVyqMzhRvG8/9z4xdg7T059QZ4UEo/9zsQcQA20
SqvpIrU77d3eU7Kt+6+H2DzhC1AoWXS8vKwrL9/UPaUkbFKcbThL9v5DB3/K4jOOBOkCexarez57
0ajTDKLY70If9yNfwWYSIjG1vuU0OdxU0EhjacVFrW80C+vbxFaLMPXyomIhvivrdDGVQFETttm8
G+v11GH7v+3iuRuO591BCLNNE7/dapMcNFWLY8y37v8ExY45gqhi3RiW/hBX+Rq3+NwpINZ5GlaY
DHkmYSdFTZZmNLzRscwkl4jcq1Id7sZyAFoQyVo3cXaVifStZyrjz2611ATkBwXT+vPSsqcnwDeO
BaooCgjSITpTzzNRUJSQwyJV4hMHM9TSjSB5wMZgbwRFy05SFunRtsRRyG2Q6QYGOrojsW6fYNLE
yB3YYdwT0AOYfLKJr2CWfzUJ3WjoNqRJffgjEipHxo5I2F2RCAT3Ks1ZmyqHOBPtMq+WeSAO7o0G
u/2mULcgaue37tHgDVThl9zrhcqPstjPXwN4mF3S6tIwnuDR+F6i+9tgwyaj4TG2QX+siJ6NWbRV
Ke+UswUmcYLWMFJaqK2vrGyXmLnXSuhboXSdMR/NoEmFbhXBBytCXBrkbh10fayH8qZsQ3J7tYHM
Y7T27Kk8MVuVMd8Wgby0gOqdHBYeiuaRRyCEsGDGK0pfFi6x8QEK6I4RcwVGx+hcyGQqNOuxteXn
CXgRDKqlMXRziToCXzCqy2evtAYwSeskmHPZxusL/MqncYoa1oax9kbDudYDKp5cJ+5s2n6MHEBI
IqyXfjXOM4Qf746Ris5Mi4ms4AQot5RYtpCgW7g4zTAQFmjHPqtxtMo7mFNkw7WgJYCkXUdEvDVu
1dy1dyNcjQVGcFTVp0PdGNjGWxvwcLOwLoE/Gmdax/c4EMdpY8wnaBLUGpBtM7gTFBjA1HTPjJXZ
UmR9eZzX6uysLBYqaPlisZ8H8+/x8RP3jAuyR+g+fvbAfHWHgK/0/xYUoWKsGpASHdMbZ19v2EqS
hTKbQMqcheC4H11adSvXb5QWNJv4Y6cGFZAndKhQpdDppgIiRfO/5Rr+HoWnccDcfeCH/p4DdSZM
1yQy8tLXBho81uWCMC5U5gbyDmCYmSQDsDwbKQAtLyAHKyuoPr8nKhy1WVvCWCpe7Q6Ho32qcxvM
Uu9n0DXU3tkeZppn6zmaTvdfiUTgJUTESVsQZOiVM5fB5CFTWwTQzFIHY849lwcIf8ycO99L+SrZ
ZpjxYrVLYfU2/T1CC9NRfRaxDFvCrGvWijgZMe9zvmvlgEZJ7ovFOQ/TQvr2AJyVpE1EGsjp5Kge
SRjL4689n5t3N4L78IHjrK/puHLQrEje4AWbBqPukoORBNcQ8blKNJECgbhOBvSAgNypH7EWOoM8
NZJHQbpYGhk44Y244rCk8HjG0oJD2jj8S/yKnciu00ojNR4uehi/nuCYnNoo0dTT+9LXjXF28WkI
z62nLaNop4j0IFfIp2YVv2G3mAnQ7yZ1CCR+7xOba7YwLFTl4gb4heufnkALH1/EPSH4ustc9hw2
5+Fy9WktKkxqZ7PJ+wmZIYswTJkPdMdXyiIIXuHYTa6HzAY7khQxN3sh0MLcorsSywaNRhgnM2s8
TZ7KHv3Q6gtcnbu/QGvu/8h4nbZT9Fne7JBsMfZENXbtSTBCI94A0Q8qp8u+a0PgxCT3yjMdJcWh
O1+dfnG8oYUe2ZD0YgSOxXq0dxWHXpNqsm/lNL7y5ffPwQ+LWV6Dzk4Z3BMYIfcPPXq8kB1qBGb3
l+vpMQGjZ/WLIOWunm+jLz4xX9wkEzXU7RozNpPQKPc48tRxw4B3VP/Kf6yoBWxkDIBpliMhtbSt
xaZ1L219QBl7SUyS6jl6q75KeKS3KwNc2L3R2SaZy5L7NSPumVkx+W4KlU8heTq3vFD8RSDmt42q
O7KeO3AXr7v78gdCU37bynJ4cwhH6X+jGpXiwnbmoiAohT/Jii4QJ1CjV6T/tnBtTDy0tu7Mkmrj
Xb8wXwqOnEFhuJurRWjWU8p5kRGTZBUbMkT+GaTNh3YGlm0lIGc5eYb5zVw0Vg6mXtXOu2VbhTCr
8hioaymmL91utg6l+jIKIQBjKA2eP3M0siKtpkwc7S7HapncEX+HrD0d1Z/lj1aqmXMCjPyktg13
1R6opFazsmjYAjlMVHfEgkEqNYJxqndW8RxkEztE9manAYsDBpNPqdLIa74oyKovlDNP9tlPteju
rk0EARdlXSKZLo6T7O/U+2fFRpJQ3vUBn3hMTiO8inJoofsEykNC4rPmrsmh48puKSKCLoHujueM
oeI+PTiqDInKtvwB12Nb4rcM5cSC5nxSWeNexQaUGgTrw1CKwBg2K7LbHxuQFswMSIJSkJkX/w5O
B/u2hxMs85hDsOysAFQdZ3B+VgArhhzYYjlPFEMCS43SVT4bkK1ZBmYchkxeCiAN2cGT817gTdE4
06fUOEWCWEpN75Ze8xKbIaMvEDzn+gmtwFp6d9k7GKRs8nIQDi9x6cncWz1ggR2IeEQOMo9yuJVF
uzTSWjSh/cY/xKiKxzc07o9yhW/1ZMU7h0U2jtj3SClGwTkh/Q0MMcvdXfUNGu0q7lk+rqAtNPMq
uAyjwofkXwnGEzgGj+P2BLPBkqkJaBvdLPF/Y2R8JyV4RzXKJltcj3Jrk/g2KZ1GEkFZOzt1ZWGf
HYj7U84yl/ZD1b674gk1xB8JBTvJZAtlp+RfL8sTqt2PaA9cDXzEroMVSzvLRLNOetz+BGQUqwmI
cv9x34gWoRY4V3HG6Gni0naoBiphXQWwhEXBhgeW+AetCmuQjOtpK8h9cFu0DMQOt3cl38JO8vol
bZ5vMbxXeS2Vmt9+AofFZBBpR1LDT+f5t5kC4PUo3e7+YYYLUEMRtjaVMddbdeW/s0kbu7m55KTS
2TKi8EB2fngEVgsb6LmjRSwp3EL0o9kA/ifCXcVYpWgik1ojuE5XzrUP3QNgOAVtoShUf1ukp3lz
SlcjCuHItOtAKCU/Dpyuz51CT82vUdlPnEOPWi3Jm1vmIu7pEA851nCudEX2U9vEV8sESiqxQnf9
CcISwXmNzu+po4qHSGXNCYnKlia6xXG9tsIADL8acZBbX+7mymLk0y0UX/c6Sl+H2fcLTVLoYUeX
Bn0qUNrIkh0Bz9Mg9lf+Vps5MjlIELXqf7o+qO7pWYn374lqPrfA3T35xBfSY5j5a884QbybRy8Z
K6QC28f+RtgEssY5tRg53lPT/nC585QZdBL7J1gjqlKcKTxGDma7ctNx2IS7auqVWGVdZuMes8GU
3R/pn4hC7OtDV8ZGsUcMmt+eTVs4zNR1MFOocRIacBpiBMeA1Cf6CN1aahrBFhh6Q+EshIAqoml4
mjyfO269Xef81nVxb8QSEkaKHYizdGEKy7zkPXmsHPcOxyTKvi2TcejWs+TrAGDxs1fJJhl8L9ji
+m98WMkIkHgVUOOVTisEarrWIIJrKacinFFPpFz48qwBhDBwOHiurL0VYZmbT8+y7zGGQUWXq9Un
jnqduxX3pwZ4yVcDkJ5wehyFhv9PwcDaQzFlXSUYGoQQ3nRsuIaM3QWEiEy+hbFSdMCv9orst0Ab
WKcu+wAMswl7uVmKWVAOZKxjHqcTpo58xeNrN5ZsvaIPETjnR3B0YWVGoo0mwvNI8yY2F9Y0BsVQ
8EF5wIqzj1ErkQjpmsCJTwT5smvYLJVTgyCP2wHdp7RZFw/M7Eu/cVuJ2F++vBjNrETKOBF7cJvz
1gIhf5HyJNQ/bLKyM+oNZ5D+uh6lyF59TWIMU+mz48H8AQXO52KGpwRnQhzDJQJ2TyZnpRqwna9o
mw2i+bhbb/00GPEomLyfEe8iHOVIfyfAKvbKbXfrphPmvlHp8Ia2FEagolJZHtlfk3CwWx3rJUr0
DGNRC+panYx8E4QJ56fgjyk8PsQi7PnaoDraNR45+K8QQrZC0njzntkq88N9/88KoRFpiroRmsLr
Hd+AK2B2VAf9qnwFjZeAPDPQCdTBswLrz7DLWUrd4C8tZ4bPUc9ODWZuMI6DTIT2+/LgZLlORPH2
LDyzHAF9ERrP9BA0wH68jty1Qbl98VkQ+0Utsn6gEORDgThB2oy3pyhuqU7lRH88/qyhskI4Z+Ja
u6oOHt6HAb9qq/ud5hvVsJJwxGNmnoH5zlc+Reg79tv1rWQRxd19sjnF9jm747b6p1n/7bs2ZBK/
zBbHZ8DGN909HqdIqVtzWG590UKJWwLXc8/68Ez5rHUJrvXZB3IGT1A3+qrWMj+aRhcDFwSsUQrs
GdqAuJ1bVmzRE75Mv2lbuo/xP7r1+R46bK6R4KAoyFmjzYw+GEgenQLxWrCs9SvdEwou5DG6UUjW
pHtEt0LbKxBoYQkzQ9KYCzErfCM9doWJicaUNJ65Yvz37XApiB3/kN4LenWJTBLiDPIV6s/FfegF
XsUERYsJ005Eoy1oG4d3I1ZdJsLKmFUBWIfPLo5K/ORRvLfYaGkyxSnbUIoUEg6Aj7Bvk2O64su2
OTuIv7C2xhrBhrgmeIVC98zAtzorY8taM94uxXJKYko2wyoZlQFLr/utuh1rVFnXdk1olJZW17km
lr2m9mKOGObSmpeKnAlGHXtYaCKjM0gxXLp8JnyiR7+ZPUToqh1UMnlTMycuLhCQbwkvqzP8fyx6
3axCxD73YaR8/RwCsxsOw8bZsvcfA/4Fs2PeFpeYdFnq4j9wduzpHVr+LwXzZ4gWAsR7ev2uE8Ep
jDh/2JeqILXiNghfZJZS5zuxzhZNosroMYnLcWr/woRMaC0AtFmcNqfwylJCPxAC5O3B7gVWS//f
c2THhskF6clRvdDg2VVDvUCKujNzblMgMzJ0tKUnsNJ94S4EztXwZ6c5N+b8QH/JdGft4s9U+v2Y
DCOpZcBTiBIviD3dO5SbOgX/knxeDrHnoIXnqQFtxx1qT7GdLpXk1VwCd6eKrUfls4oWVOQxw53z
ts44SikkR9YKsmXgqkYfl13i6OYK3lW52QKRw5JD67c8QrnsIifsL1X/gCR2isCIEPPWk7ZwFHZQ
J/98UFKQz/WJYPwtAKOX3KN+8CinunbNJJjVM6WeJPXfFdTwdwt0s5XbyV7y1KqP4lmkzBLX8ysb
u16Ge9ikEq+5GnvSWNPx7cFt37UzJGeJNo1siPLMu2IjgagskLgMRN4LGvZlhbiWNhAx1amDValZ
Y11UVwUUOZQD2jynSlCz2/aEju4oP5GsD1PnT0TkdmyNs+InPl2/8Zqa6Uq2tWHvHmobV53sixr8
EYD+7ZNPP1+H4sSAm4nK8oM/kg1qj5gxqg/UpBmw5eU6WelUA7aotsjQtSe6soVTPdIE9tfEpHPJ
KpfYHDf0FJ/tYv0kt4aJFxTl2t8c/4WfcfYlKbuMEwCsjTTeJ1o9qzK1x7QX7sO1c7sQdk47CYWc
dm/Ud6085j/CtgpXER0EkHxijFP3mT98/9BFWTfNjBfvIpK/ERKHc4mWwzyMCcxLPl3efhjLfJ51
EhGdVrUgzmFEddTZDq0Ew2KwPzvi5+NZGLVaxoSiUlf6+FMPfSYkwf3Atd6tMGfvtD77ZslySCAj
kgn6QBjg4wUTW+r1JApPcoqVKv6cCMx+HToYJ/qxZ/WitntVNHJCzCmSXB3drzr2O6dV5JbBi6cX
UnBGNmDBIbaPzyTtQ9xiGusudrUvhZZCtxyjGC149FOIT3Ot3NQ+AW7fGmf3KuSyqR78NfGBVdVL
OPlmpD5YgmJsfK8RQXTzuwj7XDyz6pk5kE1IlZqqqyobvLgDQbi7c/5ivCCqvcetrFWkbfXJ/WFO
tuKpguTccMyra825LDENUXMR+X2ckhuvx7LQs8w+y24oRooGAj/Y0BOTQrhGxa418mTdyGSUua50
B3Rm8WPgj2r+xoS0OpWfyqKwpap10fds0DLxzJLgmYoHYQlI6xIqdvHvaxQmSOxr0ajR9Xu1dyQE
QcXe3LZ4WmCsSMEzEiLqsslDmfnXvtwcBiKZe542ZObOfoSnRG6pj1/OYXGYbT7FqZJkjPKPNj1e
y+BsAOX4To20I0NGb7vbMUmYS6eta0RpNzO1JP6twOqdqV1tgIc6y8GTo7uqNocd7sQp0nfiK/TV
q3pXa3i5kAQGjLyDPGyE6I9WhS0ljXokK9UWVfyLTM0kCCwEgafaagkAIB5BBaZQ/2n3c8pH5JDv
XAxNQ726lWljKYdvYaZShQE9sRpzXuZ11UAootHI8Xla6LP/SFODX13uAHjoQH0GuM99ZNJ1oHOv
matb+V26yzjowjq+KXzliQKcnwP+kX+GfHOuP+I1agL9FydNvUhM599SVa5JxfAvkUToCq8eIt0I
I/kwGmGUggiTaCi6UnlWGyDbcO6jCfhT/GzlQ5s2mViAgEDnTLfmuRG/S9jk7Mfp8ECbxlcoZGEY
VFnQQbWepu/3Zp4iVTn9mbYgaGgZfCunV7jHrTGJvt/UK7KVTjYtoEC+6w5aaKJuwQ/Lshj4Utry
IZSt3Z0zH6VaPFd2UwJ3mCiH6vfi+v5eRQTz7ggSzk61mgGoHfS8XG0mc9rTpfUCEdPMcBVPj5W6
GCqhKnnYAGFSZ6wSuJF8L8Y9ximD0OeATVPk0V5S5H5kYw68Yd4owAhQ0wnKh8XU6mSyz4/q16qz
mSwGw26VkZILd5vWKPjIq3jhlpPGWhnkdM3M6yoG0n/2I2IMypRNKBS22+7+55s5SlEFmpKm/u/E
wxM5z/3jBMyV3a0N2y+Lme/SRuHxnRPKazoS8UlZReNMx7vfbzIGem2BSityZpXfsAR0q1KOOipV
D0vnmciBiU91Z/8S/3gWu07WwphSIaMatB0QUaZNTh1Xn1bCM+4vSCFDhcUy6SVNq43cRhjDY9Kt
RCMisB6z69/+LdQIr3UIyeq7vyirBx0sQWQqDH81hprA/q46j6B0W5XOJOUymHYHNVnjZzowoFp5
+3qjuNoOlZS93vtEcaV9JgstuGYKzGbp0P3oaz+uXdOPwnpfQRQr2vTZoygTOKp1SFIHDj1FpS6a
onnUsvMO+eDpe93hwIHkT2qak6XrV6wxMmfFK+KhIosZ+WCE+ZiQ8kFct2ze3RN83AmP1RVmgeYb
sUD2DnK2zXqgHR/y0nPkzhx5Q1wpdMrGhNdrHq4caXrLWIQ7rXakD9RbDrnjQrW3r7fPXsDpASCH
SeK7r9SML/bYH0jo+izRLziJQ3ZQ2Qwfn/bT6tPNyZTLuYvrgOMc3r6/b50GEDbHE5g05mpPM/07
w0MI1ZnbfVmoYTqDb46F2cKc4ajCjKom7ZGgpYMuiz0AuZbhvGl9FYKTrgjS2gLgnuHFTwZi+swP
JFKf5sHubfieFUgAMFaFehzzIIOlW/vOPSsLmrxgjjtMBhiWdUyA8zJnr8LuXhxNjFLCWgXa+lCh
Ua/raGvv21HIlqrcFNVjWXkeLEAwIYMRVoOtPc9M/CSMhqhXLse4Ovak0qWqD8qkKmBRXU2BgT9r
jMlFLP+TxFayChOdeZUDUhQ7QkRF57HbMRfsQqcEqMme7aG33Nth/cgtX1Co7uXNHl2+EJ9d862X
qdwOXD5ByNc6HnfVLdlNz6sd/uVaCMmzLMhJjSyU8mEaKrsPW9giKYIguxnGGdotnLcr7RB3Dde2
rUN2ns2xGkkJYHGEgdhvfYjTM47+8gki26wdlbHapkCjtrNQw12abM/n3G7PQ64m1KBfqRbr4KZH
vK7+aGMeub4+k1tmVZjokqBdfl0MEa1UN08hMuw7wMUid6OqRzZag5JLdsdPiRbJlxjnzo4QCS+G
djWWzLn7dLhPAN7cqRH2YBDs9bqwj3f3QNgm6lboGnzx8Mriu+t+l0Vpw8rQN3Zgdoih/dxBT+lq
zZLz2r+YTxzV0oZjk6gRBi+wZQ4gqYkRbTJcRK7cwki4MiWC1L8bFMn8q9fejJZMPepJMbbLcELd
VH3eUzlBZ6TpoV7O3Jnc833NQ2vFyttrEvfgsZCigs7fF7uuyETN8kA8DHLQGsOAK+AfR6WDiTh/
oNI7Jmh9rzs5EDGDCTQ7H7eoUN72SKRDgqjnEhZ0SvRiSMWmguxLi0U5uAiqA+59jx8jEwyz+8VX
iUpW/Pf59S70ijJBdoRmelTamGRoqqGVz079wotPQkuH0waJqwRmnrYUgKmXlg8MnfL/zgJiXFKf
OoKEhm82yMiow49NelXQlLrLhly6lvavaqkyEWWJF4+zLrafHd806fapiZPxA0HE7XmmoZ400B2i
UBGQsl9tfnCSZPLoUjElpguaSfcoMi8uX82dXZd7503wXgsx1zYaHCaNQLJ74vxNlOmUrM/lNkcA
VNauV+ZRSWNFMWJzTyRkTuo9ghPrINXlGDDUCjyUmDDLLdr/ym4nHZqyEuM0C3ipRfTz2ey5kvtl
qNQpO1Gn5HMQkCwGpEzFvJusFdO1RSndopW3ZiQTCv/4GI0ljg+2xEEOthZ6yTQ/ahIPUJ0I/MOG
P9bxLlKqh/cDtramfKJXJpWZCsuuPP7Yg6PNiP0vA5JbObxQugN2EiyfRAp7RUlFCKo+3UyZnWUs
yKHVA/AERGhzUIIz1CKFOW4gIqXBKg+USG8dHNo++nWgZfuEcNBnS4Ht+Se3j34wqIptze2Nau9m
KTwgodkEptNfpPOndxGSGu7l4QMtg9mzl85tamXgNEC0DKtANKZ+z8qxT+X/EnmP2rrxb5AX+zwo
9eC0tiwGiefUvczoriTzaKUz1iGhN2tPSWWsygk7JCp4vLcqBmCkOj8amKNzgyC/SnYXvquf22nd
niqlQNW3+vR+Qk6yt9Ur+jJwuJTf90x0fD6Na7p3NSWqAzrI85i/ofT1mlf8E+w6Mp9SaOrk9D4I
KOVGGIyf7NIb6bukOuoipVKzQAIVTtjTlO242WOBeoPYxjo1jwPbsOKugvz1xx4uHEisjYRJJUYp
bRQZJKhavQMDd0PrMzrTesPigJoOqgwB7HS8WkGtGFQCXm2966ihQhgUdq5fb1tIRZRdEJ96CspP
Q8TPEHWcLfGu2wnhKGqEuH4TQvVp2lRt9+boZ6Aixx80TXiXS3jax3AeJ6IC8YrhwShwpbHIHK+0
/8jyDv6aUZhEjd9w1RAshDb0Lm1DCSHSvrx4ofFKbW7iOQJd6jtOX7tLaN1hkpCXPicTc2nnd5gk
Y58/xHZNmg2BX4fdxSW3i57lnfdVw+MbA1bfBaB5OKC+1j1NDRcP75E580PNzsrjsI574rp0Uq7a
Pg9i0rKGy8BHpcKa0kh8vWnGJYNX4V5fwh5RRopF5HjBgb8/24P3xDP8rloBmkYUhoD1qM6EPGEn
bS8EwLorLE0y72um//n2S15WpWpHuRMTzp2aLI8a1mnvhFwR6A3C1ZXu6FPWe44TzJ1DCJnh1NuB
xtHRKu27wtkkNAcRcu/hnsaMxMnVe1LpG8az25iuAyJlUksIye2C4sTZDKUEetUQ95C+Ddj6B2N5
Y6MJ1T0ZXVbx8knwZ0g3HNj1tJ08bkhLI4wwszg25h6KnpdwtgYLfYVSt8zMv42GtPqOOgVzCXpt
KnJYGUgMdK5D8PoD8oykHGjVyte9TyA19UCNuYXdgVt2HRYlwMLBADV/5CQxtGC8QCfuQZ3GG+Yp
NhLFZ0DUWs4/JPWxOZ/C+Q/2cyhd2fXRj4gM5pAuclpGyxKYlD+mrnCD9sh0lbNVoHBLo73gt6Bf
xjwGcKAgKJxl+tFMTIlyyykGqmtV9yhlyDdrWz1ZfOKIcrohJBbwoQWkeQuhsChdLMZrr5l2GTJl
j3dEbHqDUcsGowac42bNpsp9Vb3t8Mtts4UbAhRfbCHK04AY8NgYvcIyWr7yK71reByT4LRYMX7B
Lw2btLHVHdn1JMwI+vLpCOOI45NAXxrbwA4mZJJ1wc5jRWE9utwZNq4TLRa4ol5QO4yEMw3CsBRN
O9HFdQaGYNOC95WmNkzvAMCS92U7KeDYCdxvOuHFTJR3gs7c1BLrSfc+my/ASpO7cX9ZKGDQ0mw3
D2cXfh4lrc9iVGfzjbWaWbT8/tP6fFE9xIosYci3e8nmY1JEqNBSAswYRIytZIwUUEidCu0DkFcW
czKx2ccuHNS+fHFWqf8QvJkImCiFbMlGAUNIuRzEa13cgohmr/YBSLso5F+cN3nGia87r+ivUemt
zk307rRFPZnaTDZQYo3rOrZCxAGbGONYk1VJasTYmjyEd/fC6sOgcaAWlJdQFGDoycR8fHYDPWJs
/rs6cYVk0zROwMDbw44ksF1z2KC3973kQpkvq7NgDqNV3XnMvVImUQWQ9Cne0+q3beFNriJpQrcK
75ydK+2ioN6WOxHCqPXC45Gxt+Zrw5OEdOrUvFmeu6eow5e/T22bRzbO/e8qfb5YLZHd3AX9LHIa
9NM9067VOuwV27QlshFE1e59Cf6dNkyvELS/JkKLyrEl/LcqSlNaBdJyMUSSE03XrucGfQOvIYdG
hfco9bRLFJaUbUASDsgsljhF9+u7o0o2PpyR+P/0rVOh0qkBcYdwh7BN7R9bGgxeywLlymNayrks
KP/CuKuJMngxI06ULmRGko2/Pxndx5FUrKbV9HqzmnXl6b4gBla84AZM0Q0Pex1ZlNV4VflFPkEf
3Xh+xiQMMqsVE2BQ3KE03TJE/amMSROfoB8Npj9xthmxpoz3sIAI6Z7ckwoXi1UbgXcy+6r7sxw7
1QZ8rez2N1J5DZMPD6FRv3Viq52vHz/J39F4TCJVA24EZEncCYsqV7p+ChP6tj0XVTuPi3cBffNH
J015/GZ3PKD1P+mVoxJyS0UJE7PDK+GFhq15I8eph474FQ0XLDPN4vttXS0uiEGaHvLTgXOrOhhu
cTCgBdkewJTu3i4ghQiIC7PlNJgsKvNLJQ4aWG9OE4KHfOc2E3tGBOVV7THlCUDljmlxB/lFjIUI
B4gG8swdQb7YRjADneBdzLddnkApay9PNuSQauCNhZjvzAQyF42Vm2KEWbwsfk91aqg7VniN/n7T
5i/cOcPu18dKGl/bNKVepRtZGf6+/z9kdhubTW56jdHgMo8DZRlgnUKqNrA+xfNDABklcri4TX8h
es8KuXI1KPRS8E6DPP5D0Kc6Whm7rDbfReur9P7hgmOh1YMWA++Zyl/EgnSk42EFNJh08USUexWG
+NZa+ULA3RI4AQPqz2nGsasPG3vKhbRN6ZEj8hYHvsIfytC5tgp+DKiLx9vQdBUfoxF9vMjRAGgO
nqekSmEPJmg+3EyGfc2P/JKwBOe5V5tZi1ozn8vBrltDqW7HQ6PHlOK+6Q/fXHq8U/H+1btZrYQB
Ea0x/muyiA8I5Wdc9UWkHI+/4cjdW2TlFtELGSGhHVGy9bC10PH9UJ98hTmgkPhTgmUURVr47T90
H5L6ijBifCDe7lJTMVcZc7PZ6wKRemII/mdshDoGTm2lWPcw8Ad09gISpwJljQD5xTe4rUJBkIof
wLp+8KpHpwpqI1oRZ0EVLeX1PwBTADr2dx0I+tjbdL4pv+5ieyNU6bsb02SannBG+WVQfO+Ve/Gt
Ur55L9pqjNQX2sJ9plpernHrxrJ2ahLoaQlgZ/t+sRnN2nqir3ML05nkMWfyKkZCnJw8ZWJOWSui
9jWjYawn7Hkr628PEN5g+DtnzrByBqqL7wqsEIwdG/iL/vaJKrAn6Pl24o4X0Lq02ZUwwKkc5muF
q5CjRgGbLdhsJPWJIwa3D4tpgxN/cKcoV/H5QlLeaD+EXiODM8HgOcvjcTfBYETU5jN5vpSpJTES
XyEbfQKmp8isLRZBtf2Yz6IJf5vGi3afRh4u3l9jizN/i8I7FZzIC18w9vOhvOhPd+hwTyMhklGD
PFCKXTlakG5uJJGHPxMzNZgZK/sZlpiSGMz+yxKP2qr8cBZ7oacIddrbdQLinTGznzhST+2CCRXg
LS4+rocZyTB7dEH2oTbMkbn0wMOrS9YCSi+l7wXbF43/iWbg/rfA7sK8jaCtElQ6y/xAh7HoHUXm
1DwruMRz6ptjcPL+EKryoSUJQ0IziDuCStt7vA0wr+sMH4XBdUJFt44BtWe9XYUCXnakqSkNUEBY
XQA66FxOFoD8/6hd/SESPd1dZoIacYvo+z3DgBcA8/nXpYotA9F+7NyqW63lWvpfI+LqhYhLJfIr
AVcAD+3tuh3S30KCdwqvz6zxFR++GAvUUmeaJneJCTpP0JB7RAROtH5yXrJqNpkbl9Zo+eFWmuJ4
zEn4F9GFOckfSQ5imz0UuhTsI8W2rRs3uzUkzEn8RfPHZAPSL6EQxg7aDqvvnKUHTEOyGrG85J0p
Qo7Ugi5KIaGVHJOEVGmEDXlDJ6tpVVJhJ4lIRu/9WIp3V67nTzZdl42s3LghYOBHWo9nz5VkMxdX
lK3cqTA9VIF099gY5uEn6q0z7X1CMtuzkdnunlHB+A4fRMWHf/Rj4PGE3SIEqi2ekXwvbPBTui4T
ml5WdmdG+q9jejzExAa3Q1lQj7eMHJFUDyW8vRfpT8YT8WKtLB5BxPdoA9UUspFrhdOPE/22HqM2
rs07K8Mur7CQbhINOnngk9AghImQPXeTKQIdBXkHgSqVsHOE3Ub4vjYfE2wQ06OSyoJeTFcy9Bwo
LR8S67fRKZSEcfMoU/0tlUkCmtwKQpuO2DD6wwu09Y4xzPtVClZrZlqP6OTwRlYJdshLrn5E24BR
rzbZoXxptxixj1XYviu14yTFozemhLSbfDTQzC+tsfswG09kuxiCrqbCukEsKjqVWjZq+0J3F+qp
ZooJH2lR/HTX91ZNPjfzXWkAeCv8x45KpHJ6QvmuW8fcZ2WjCaGkBrw+czeWINBXEng8NQGYHzGY
JR+ydc2NpHFJyczsqY9G1M6PymI0ltjfsxs5MepZldWDdNM+AloqZ+a2N12f1AkdWdXrz3A9WSSb
fu4swnKX5Jm2U17xVZxdaQLY49wm/QcMPSv1fQN/Qwsl3GVwCLzYerlVMxukSdjwwabeueE1lIsi
LgfsfIcNIRsT1Hx6dX6UWGvIX/MT+AaITa+A7EYOGunw7YOofc7fisbvFOg583VkSOE49hhZq8Ir
HKgy0CyvCX6Y5DJtI/UJnoJaAhZNT/Ln0/qjqUY/CR79FjD9bKSqj3hirzln61zj74And7mieE7W
uGHMK+cbdlBPT9k6jsxZDqWsJiRCiJx74ljYISNbInZJwVuvGIJgXPmJw3Gau0j3eo2D04mFFwNa
RE6yo8aI2gQG1RCSHKQwniB2BzRJxl1Fsl3oqCZ+5gaGsOVdD/XVavobF+xXoezfO1fymdKkuh6M
L8a04V4Fekq/xeoF/42ggba0iJcNJt1MhT2KRJDj8qFsK0YRq39ljhSWSCVoUYjvOq51q/0clKtM
4HFlJM90ObFaiZjm16qBFu0141PS2Ies2oInIqK2jNAfyE41UFT/C4Yv3L0zs1x2PRQVeKYP5R/D
LaPShEGqVDshYpJA+SNlFoH292FA1SJGxDAXIk1GnW2HouxjrQCrb4/3WbJ24DmKmxGS5Hocnc0J
TyZA1B5HNkOcnsoiOA45BWQ2v/4svrUgTsHUnkNioJMDN+6jpdaz0tKCt0VoNSpZnPqE6qibdGTx
g3YiGtbp6PgIHs8c5DBbmzhuaurvTRxoyqoJVPSv2t4KPuE/P0MfcH1Y+r265kstN/9cvtPnUuWB
87Bo8TuT7wr7d5divgbwhjMMOyH2hSzis7IHIbqhdeYuewPRNB8HyLyBcSP8metBJ77wNr/Odlmh
Qbfyq4nzDOiYQowMFeVbfB6X6EiICvtZFwZa/iTUMzJEYsnZf2xr2EbnUP8eEABFnHdBhglbSLGA
QKhmGwUu+LnXG4wtDP61OWeP0p7Kalet3WE67OgFit1XadgfZnLRYj/z4OcCFcqxDbcY3hhcf/D+
q6xU00NvwtZODBjh2KJgbVPHlbjnmu0TUYTvR3NC8FdjTWvGGVYr4RtCUtd2rUGDj5dL0s8wYSzj
RFVRHrNqAmRclluLto5mEYG4XWPiAmY76GMILiKp1ShOkiH+mqr1pIOTiT3+02ISVRQckwJ7Una/
hyTfARH2ZBe+GRbuQJdEDoaGKUasyYcYqRdC6TdYIx/Lfj3t9z9miRcC/WhStCa5KXfSo4yRmVxv
C4MHaf5YtrrrYmZMgofKn2OhQYPGGtDSy11L1Nj/hjGIYsOirG3t1Jw6DqnvlKZqtK1W9aBR5lO1
L4S1jM9ygqKf3YtIo3jJs9Rvu6R4L1Gpzi+VRwu5GRom/uEugVFMwdqLjXr1SNSHAx24t35GcK1T
CQTfU1kOChXVkS1XDOu6p4fmoZnW0yd6W6cDaioXQD6l24dcOFAu7LI2K91W02RYW9AJlNp+XDFV
otsmFyb7Lf2dhyFQt5CwoNfzoxZVaRAgqmI+zuQ4Ma1KZQvN7cRPRiFA8vJ/ywX1+aDQQmX+KORO
gDinnb8+38oPEKEIb0YJrh7aaY5vnEwaGsheN9uEQEOJ4WZ/zegVWQcqupGfGT8AI8wydifqkmqw
1Uksuguopf+iCIPwRo3bs6b+p+FxVn0PjLrJCEsIE6Ut1w7xhCYn9YsBzDvFv/Zhod/yGKZhzXlZ
HRftX9OmGT4wWKw8xDSOfXys1Wz4xuN4fWU59YTLOjgYU95VJc8aTHEtqlmwa8XDQscs4x3Gtqov
9bgu8n+4p2F/ZXm9LxiB5+ZTa9agK2cUXLvuopWoQl7fHumw+x7LADhXyvs2VP4HYdqzSGjw7TqW
wREIEamOS60SkL5E81AsTY43RtJkz9cubeRUstkRheqgPHlOLGKiBNh8QzUQ1QVKZhs0gzM7qANF
GiKOr4DSnEPkZOKfdH4vlnS2TqQH/DEmi/HjLtPS7hvvLMOeBU93qxrTDiJrICJP/T60xkDjpRQY
+xAzpSCGz9iECNYuPrsak3m/tT5Riw1w0X4QBHmKBSoV4ueoSdhmuCVKqi1thz4nZY1v7p7ux6NI
+FwaNQ1uUDyFFYzfrVOpZqU7+5dejK+F2eWzPQF5Zb6kFGl987k2MXMrs28BAReCrtEHFxdUIoor
Mf1I+rIrj/rjv4oCMS45XKrsecl3WRA+ipYCfSe1w+a64x1batSkW43h9yt0R2jnBXDmKBGOXl7h
CoCzvNerrzwUAyrSCIPajKLcgUz13mQhl4WqgGedMY2k/qilCQK26mDkla+6lM7MGCuROTYDcsQD
rvJMSZO/81ItMkYHykExlTjVpc418H6CkXDUkkwWbkFpI03+KXgl40O1jy3xMpdMf7wOBPjKcTqY
94GfHTaKBNbNDSySpdPDYjoyReymBAjp+AyFoXiKe1EQoIwRyk303H0aTEu5naSCi2uGoWvPwLLE
8UeJuEdquV9VXgdko+1UPyeWcJHzlqtMM9IpGzMHjngBlOpmvgXVngAcXPJXhY2/uH4sTcNFAv8G
8UpNFcclV8tN09ShkXE7q8HmSeYsl1nM77g15kKcPe4X9rad4hAEcsoR8fQHd22x4axCnfu3/cHk
OAaNOKTMkuWWncwCfXXjsP12ucwkxaKe0pr06fSan+KXxvPtqSEz9oGzej36TpHmx3HorCsTtcHk
5a/RCqn1jtEpg65uvqZUs00D6AWBojiVDnF+O5Jeff2QMmnbY73Zmdftbpb602yHnpfgrdq03V3z
livbRD2JZlPt9wv93pdaeVCUdf4bQfAKqrcdUlfZB5Sezum6jfhgzjGR2HUUUBw7fYhEORsGPWcg
pp5KyXBW7l1Zyh4nNO463iuPZSxiTGR00UQbM4IgFjD8OycWBiBYZ2oElAgbIPzKCSEeSE3ydCxo
Fj0OT2qzgaEWLhVRrAwsweA6HATHfkxZpOxoZzhwvOwQ9d6oIZgiMg9ApKmTRN9RJe2o28wnK/qZ
ReCzlDZCb+ltLD4A/7uuCx2cGG6VM9fcdeQmyzHEfA9h6X+KLzwURjZ6mHyd4iSr1vWxrbdQgH+1
5gk2Q0cWt9uMV7pB3ygC739Chcfm4GfZjDQ3/D3omJ1HDFw7hvv8Si5LMqQGYDuV6yOU0QqwARIo
RcXmNT8GDsH3gKsOYKsMuvMdJfkvWA5N4ShOSur69snz7MnnPgcrnNPGR6ry5IUd9c5EzndmIOzK
6FQYnOavx8ZKXIVOUHsWUwBVXownaOyIs48ytX+eUubqpvQcx9QaCHYg6Uph2vyvd4xDMEyuCp/G
PNCpvGFFK3hreEtd31XG9oP9UfrJQ0miVqaLnRxaJh62ZWqwR1pSPQQb+GtgZErkcojPi+V2YmNy
eBYXTW6umtaMx7ceXzHxeLSQRE7N9sSqdTW9mLqcaoK9nPOGI62JWEVZFCmooeJ9TyqDy3AKRFhg
Y6bstrpGr92GBKWP4rYi9ONv7n/PCAF0bvwqQQ955ABRRvaWLEogwb1zl+QRMcsxxwRw9mXgXAfE
q31XMzppyYwh+ASlw3MnKpAmqm1lJPfdkuESmcqE8c8gw+RO3Yz0S6HfcZ4wEZSP0jp07VtF4hW6
5iK+ZJtB9WCTsMF7hMuox/hUYJ2mI/5YGqNlzZhRnlkEzkfxwoIabMkWqQGeEgP7NrpFRvT6eB9a
m+/RucPVvg9bFTTvBquwH0UTz/2saulEUGcQqsNR79aMvcjY7a7U85h01ZPqJzsp2R8NwATluREq
/+1qi/ZGum+M94G3Cqphpn+8xMGBEBkyW3MIx4ynrtnuZep/vkNFritHDbjk7Unl7WxL6MqhtGC2
S98qnwBmi3puVhPtsaScLc8h1s5cid0HFZlvnuB2pNfN9xCcbSu4e3CvhXVH17lhr/4MOjhXb5vL
bSLGDv9P6mVWo6tQwfAeha36yVyhMrh52AVdTV93HxChYlEIVlez3gq466DruxfTk6TK3JBuyuwP
1sAMYsatmw+Z8dS1B1ZUbDqWytYu7eVfzUVELNO78LslKBx07Vss2B7x9AkfqqFeKEFcYgVEY1Rv
o1JptmKt+NwX9ODh6U0NCPJ1BXLHgM4B8g/sZcNXEGRVc52QQojV0iCYAI8Xp6LUtL/+AiuQxuZc
IHoHxPDWy7mk7r+reaX5b7Yc6fjItim4ZVokQ8A8VILgB89O8ITgNYnMiOL1C2iz1xB+Rqzp+MmG
Gq8yvLEXJv7Pu3tzZ54QK0FUHHkcjgSg0/oyWnOFIsCOgLP7AfJyQN40bjpHvFBKq9aXuv1nWFLH
8R1aotX/I5g+9bALkeHWdzOhsx+FVLrin1y0ebzq/z34+eCVlruY+CfGa6q9hkcXc5IhMxsrT1WQ
g/R4LBF+nM9+2VJwQFLOXyuUOrvhw7dk+CTYFJ/OmCeG/7qUN5mApZtjzE/zAsQ6TA1psqm9O45/
UDsfH4iO3JKiRJiiWbO4zKiyFoHcgYJrX+GN00Txl+za4Jl8FSrX30gDynZZMENgUGDFbHCwEV6N
waMID7tuDSufQcea98YW7JWK6gp67CB8U6ImDWLMW2b0UL9xd6ApD92fvUdfWrzvtf44iRnTyfv9
+4vism1KL4YVbLo9bNDwo7IbSRDWQ22+r7J54Not6AgbzpSfJ/DWqsKSEpbprS+dZc7CAGiEzyUc
RfRNG5hZomXg5OBCk9E4oqvKngD+4W0ZJCdlZku1I9z0m/PaR63zeLrlhsSnsgGgm5+h2VzCtM6e
oYiyo7J8RiUNGmrKHw3l0CSyFTAesSkmeS9CC7P+cLCvqLl29gSSlEprijuBA/PG9dosWwdrArVQ
ENMgZxUNL/4N4qeUFBQt7MIMx47rp1dEKcEPu0+Cq5npWK8GYORAjfNaugN0VUG048IRHwPfvjGZ
JNYx+Eqy4YkzoPriDTqmG87emj42DiTxaa/gLN6fFAnUJVXJvNkL9ThrWTqvnWq0ShRI3wDMXNjY
GFW4IvekHP/ctGV+ZETxix/ycuZmDAWKL2YbyyWHEO6kb4zEAr+SWd7+6TP6t4v2xaLbThyZMxiM
OfLD2zPKQ1KrRfUCACi/VEB1kj5yj45HPnzMGsFEXYGBJkQrOWBarrABIFpFO7gQc4SJngbd4Rdq
ATMoP5eSTeeShyvuVx/YzRuIjPcIPlwK58etMbfA4iknRkvwQo7e9IQmKsHvcRByAC2HKjr27St5
n55bWNs16/xKRszxGHngg4sIrJfI0qNttVqx3I3w7qU2VHLWkNTWHi6hUNDFWA8c9cINkNwu2tMY
jPzkUuVixIV4ElNl7iwdeY/5FtqfsctY1YDHmDFMJ1Xp8burhIQ70cgd/AneMit7EZ0hF0YqJOPV
Zfd/Infz7O2YcPgK7DATMDvLrkvMb/dtq4Uav6AgY+Li7eE1ChUafMZ5ecpCWDtQG037yHHcq/+n
KnfWupI1KQt7ulOvhm/5OQFcJ/H4gyiFFmn3/yxxbh1M5NiYlNEDjsqO6rE+/RdH8bBYn3Kq65l9
To4Pgj4POQvf/sLnMQSXXnnYI/+JBePXS4vFeKYKAC2y+fHCNUS5yHmyhMm6sy+pa6pfG4W10kxG
8IESbuo/CH4RV6tgOkhgS6hf/+7ZF99QA//wHJ0Rs3V/m9DXN/nsy8L4CnQ6AMC2rcQWHgwT042/
bJp0CfUjD3EaCrFuUFFTgWrOXWnwb0qAsglVsO6+KI2VJACyummNGo6J7ibNTHwrmHSny0ogIjr8
55qSZStgFn5uVm8fdJVSRwAtR5xMzQjOwbs9S3m+5BKxMzlDAeBgyBPJWkHpb924ETNPtdqbZx70
uYpRcw4+Z+hRqTCs2mtIcc2kTt3i2/qG2YFkZ/SKQ28+WhwR0NRtau+R6EneJCNdFZY68kP44AAz
w0jd0mPOw3z4MWjJXfbOPHJYqOa0S7s70Mz26JnOVYA95mDUHs0Oa/9+jfD/yo4Sk7SmmJv1QNX9
CcsoYVvEQvD/AnkdWfX6hVUWt7Qup+VC+gnakpUfSjdVcEMYezHeZnl7oFGwutqNQKW5aRL23tSk
Y9ftzTKrq8G4v4Br22E8vyaowBhd1xgdES8yjJoRYBmIjCwZ/qlshNNpGXxUl1FiGsNwx3I8ZFHE
4Ib6gn6O8/ElvQfE1K8HXjH6jckiCTUV7YEJElXolwYs9g8V9iHnE9/pRhaBi5i4lz8a95ZMPaNm
K7hMAFWaB9TLx2voSlZwy1roVrpxLNte9l8ZLOpw5+18hC10EDtevUlWnhfkpmRp8Im9sH51ZceQ
Yg1p9E2btEbhFBHv8v+8f60SMTT8Jkx8g/9vPC4cPy02GwRb9/+kJ4LtTRiMgcy+cj2y+/2Jci4w
sEF0eQvsU4v5Rp5m4WoMD3AzO9GVtH/caAJbIURxR9ALvi9Uf0xMTjXAuw9ZfCggKXmk3K6LG8UZ
biKwr3k6wig6oc1vNm5IdTZ5w/iJTfjk83WdJLIzQDHLetkZvglG/kGKTkGS4oF1V7GPFO4X5SJK
gNj5YS+Tdo1eFWN6RQt4VM1HFXsb1pOmEejqqLJ6gJtY4kFoYMNrzj+YowOHGNhw2evQwhX06CiZ
Og03afD6UqU9aUI57WSaNT5uPZJw87fr0mVNO/sU1C7dxoLYseX4tu9oC2gdHOpPWLnNhBMYZTNa
tXlev62s2SjlxEmbcQ5HqG5pfCkfPWcd/ZNutNLjS+i/CmD+TZtolqWURt3GN6sge3cDgoTymZcs
8GZSJVgxzcqbdWq6TxAEuGeGX0wSL07jDUi8VGvsFA6VEG5OWayhdMsyV2DzRK1nbQLESYWyAw1u
8t15U8hvDsF08zUcOUdaZHUEz4R/HjltkdNS9DJw3VRaV69FB3TytsXGRbdq6CzfCT9PTbZpVUkk
dc2M+QH3wHbPQ/urpINIBIHvtZfu1xBXqdi/idfkxOE2aeMbcJ5vKStdmQ5Gli3FWw6N/i9/uO7z
hV0D6cBAXt37uSnhhBfTCfPkHIgm/N6KTBW0ryFyb8uWJKBolcZqYSJVvbfTWCvRxPdC9IkzruW6
t2fd7t8m70Owm1D0nnSBZgka9UDgcfkUhhQka/r7cVQVSTNjw/6wf08MrcrU92v7v4q/jNPq4WzD
PPXzze21fEZnxAxAgDII1/F5u3m0JV+zcLAH7z/YqZNyYK0kL2sIMgUm86nhVuoFj2eo6aj6K0sM
U2KyWHURmtDmw1NoneV1uq43NYrVEF4sZyMTx+lRbr++nuhWwBe3RShKlmyZNYEWjXHPI5TS1Mig
8OpPxDT+7fCk1bJUgsfA3NexiwkfEBM2sIVNvR7EJ2NnFvjRTmYL2NjZvAKPDPEi2Z0weGIwUmXs
9ZJsYf+KjK4U78PgJE9iuVyNxH/sWOjiPvtiRuuoXuCJhKt0F44xcYJsJj9IgQOrCzfLtETkKJVI
/ifzrAk2QM+h6UMOnmMHNIXNYkQx0JYN6uk1vbcorwbEvdO46WllIMkqqno9gkZyZg/oyvlUC1HS
oSCDeM7odgHuDhSCK+HFe8M8T9JdCqr4pX2h/8aOhgH4Xlg0v/tH+Ihh0/zsYnBaDYpL90cUEf5M
9biHEegZ3BF0VBogPVsfDdzg2E3ZT2373CNOxPI8r2wKavaw4ui5TwbUJJgoqGUzwnxLDLYEy/gc
pWU4gLZ3c08LZj3zxaI4sZ8k6iA7neMBluWv54Dh6Y+5hPF12f8whqkSWLw6yKGnaxR3aDNL35SL
qN4/PFqKKgLEgwa18iqJ6LiXad5zNsvIaYH7jFO0W8Gag1WAcpCoLkUl6+DRNKv4mD5ZXQa+wGs5
yL5VCesi/8+31E73+zLkyIobOWI9hIDfElpNUDEcazn86E1zD50QE4SYOQEAHb1Z09quiRb7A47V
nEuJfQ7HsIze9N4kt4rpkdDPZrpSQ/0z4OTHDdN+7BnWSKllBMMS9NnevpB4vt7U7Axj09bvpJuv
QP/WprmG2hb70QaCVy4i90b786tMC/qtg3c9QFN/5wDxhnf6bby449ioeO3HN4Grtjm3vOBmbvaD
RgpgOoh2gFJg0VWN35JGxgdpbSD7UkkYoVKBNV+BPAzsSm4l4PA23oAyaqyuQTkaMsjl/2FP+YDM
BMyj7xz0tBRIyhHxcFS/rDdfGm7kxSk1giOxgFuSqhsVUMXi4AG+9+fIEkeKFuSq3AYSgOm0w7fz
AjRboq2aCFb8vYZvNpG0k/L5slClvtxRkoHln/yLW/Ot38fuWb+7ag5HQrP4LbxBEG9JL/hn+qYi
PruCORP8QKHSfe4huuZN2qQXbWd8mxxgFWBxQI0wdn42/Kr3qK613v+2ZvlEPXKyH9fNd2G1fHA1
zOlkvPiwUwvoKbSmIkujPv1VAO8BAocRTSU0S2ETdLqns68GKenmsTHeULWWglhnKW1jxShO7216
9GOx7bZTY0SUdF1k71IxnfhHLEcoo0ETInY/RD9+Wm2BgTpb+3g4w0lNrBLwuIJRwePT6E/lebYK
uFGQtuYIUe7MMYW9uPctMH5cY7JOT5ttTFNa2TODSl5FvX0w0moe8++8Ipa+pdKBsV9/Yl7tkU1W
O5oFPYeLSdeIPfeU1svtL4evAZ05kjLL8aLXkW79bpgkug8Y8PxUY0nMtz8vjCvzN5ep7tJ7Nol5
ODxThl1xW/duZox73ijVKCcle9at/H53yesA8W4rlLxlNIsH6S2QVJcHRynOq+Sk7xUq+gdRmnj8
Asz9F4cd1VdG+V+86JZTBFBxmZMwHovu6vQkg87Tsuy7sRzvjadbPxWdiY7VM/UmyrpEfPDVcGlF
5oGQiabKlxkp9jz8TL7/0mtL+DdzyRo8h/biIWZSDhl0UKyQsEUD7DFsvFOawgkf/VJR9GdnJV2M
09t1bMD4AMvH/mbzUOxl+4dcp2qzq1LtNDTLYQjIcBngObuiGwYt1bsyWiZ+J1KSYALdx3n6zl5b
IfodWdIR9+a2eXB/OxQzcYyFOucVB2m0F9Gho4vVdGIuNNSJbRvUbnj5axjo7Fv6O3BmJO1GJtav
bjL3ULyaB0M12zxB2Y9iArddw32mD2BO2d1uT8w+sPi9+IA/tu0FiuV5dmnnWZwLS15oDgnsDsb+
o6p4aYrgtqBZnDQ33OoBIZKVs5fA4fUuD4lrvG8BuVNbWAHsyDy0/5AYV/4zUDK+eJsNSLL6PVjq
MFN6motWNT5kQdklaMl4yxCa4JUILHBYVOy8litvkLUNuOS1AzE1PkUssVlGVrX7f9oWjgWzEmsk
vNSTC2B7UQeKlw6qL6nw8dvDx/BQxaocKX2oqqkzLhyv5dB8V7RRJlBSfEOdAF8CCF6ePqssaqU/
LlXetntJnaA/pTDERvktClwnzuzXaY3UoiibENLG+HRyInSdsw6j1jark46AazH+HOgQLJ5BaX4b
87ngHjp2wO3h/zOmgvYXkpmweR6uYaOeg9o59gzDejMS9dyUTeKLw/POx6zW7gRvsVpCZdGSfOU+
bqxGePyetCj1/dE6W6huB7t5XOlozSeFCQB57M4tLtdM52Z0gHTb37n7qK0iagl6aaicY7IoPkKf
8av/tfMdYHY+pn7zOSwX0/UVTDKCCySwcsRFbIolvFHkKb7LeFrjm386cwSO0tZm1DXesvSk6k9O
rH1N0mIrwN2tAqt1s0zyVl7f3DIA7dlhtkP3ru+IfJ8vDjHL5RKHRdLSkPpPomAg1vGeqe7LPdX7
rn2Vr/NHGHoqq6wGYUlGNhxsi3sAvnJ+VKBRy9JxVXmcglDapAGzA05oiSE+vFM3BgWUo1mCEvDM
+v3+hXGtEm3cntBJKUY+N/0st/On3zAo7Yq8p2vlJZFloZA77P8rZ9RMhb6lqoslmdOhOxB2HPc9
dDTUo3nhrPLFYbW5zEDZ6kVzjbsuSvhYX3ibefmh77JYo3VU8pfXVSqBLOpbVPC7wnTEvloEf00D
ZO27porU6dq4HwKm7x55zxH1JgIGxZlcC175lF7cl8FI2jE4cjS5Rn/wj8j1mwcMH1w9fAodIH4T
0lcnTtjMRcp4K69TghhH9r0UhdgJTPZM7QffjL1yun38NkEEWfVfaDPg4Ugds7XxAjr4Eqme46dX
BZ50pUmJIb+uJuFhTPf0Rztkv7WJJLW6QH4jBMbnPvdfSjtG55UKW0BUA1yrTh9OdlPj/lMETs88
bqmEWVgLO+nx6DYQLslE0iVfOEKRjJ5qgSkH0+FbLeo3YJ62Z5uiQA0UnJxbrd9lyDkvvwySq2qR
cdyPffr5+LxFjfOliwn/8deOThbYLuRs1MXKwAaB98c1TgHyUc8hgbsQ3LXETpVLCDJfwVbaeouu
KNUQPmJtOpSr3pRGcW6Wf1jGX72fBdvAFMSNI8WIeTUpeCW7QQIECmnY5I9t/57+K0mbP4YhIo7z
zb5JfqtBcLBap08+kMRBFo58SS54swDmelae/lWQT4apgsa0oPj2YleI07cjP0KYiMZ3+bIy7hl8
fts2wJj3ZEVd6NTtDid/mQdIPXQI80h7S5KmVPHU1uraD+B8Wll+UYxchZL0sUyOF38ySOGKr+Ij
Amlh098G5HcYm1O2flkOsbS32fqOIp8sH8mvIF8xtd/CZE+Q5bTwWv16+2OXLm+bHxSSacd8GoaP
SsSs3xzj7sS09xqqLZ/5+LsvpEQxP2VkakG2isfoPj+q6QI2yUzK2WY2e+HnWyKRZwpm+fHjSC17
IcrnhpJEQaRZbRhwGo5SzxoY6AAe7V2LUgYBXoA46xDK7Gxb7N/b4ZG6sGlWjyJhQ9eupXi2EWq4
XTvubSLZspHPYOZ4O4Otd0zTbzD0idv/q1KoneF6c+L2tq0TuB2VlZcYh9HeZEroSY9rHXW5GVp0
msoNFXng6OGD1BFSGZsr2/ka8zc6Zjk3bsM+cputcLzcE+ANEmBw20li+pk1pKrzVDyo1E8y+NB5
Ycxbh5pDNkOfdzr7d00SC3EcMAf/MUHEyg/Kp3CI99xiK5T2tbqcBgygxlJFYbH6mhQlZJUkapYR
9O5Ya+FSRMY/kB4EhW/+DqnIy4i/i0iIxnFu5tLiS+ss6SlKCOqGwsbGTP2zXgmfvJLjXKd1zlzO
GvkDqi+ihTocEpJTFYf+BVgvc/yUrDR3LeG1Buv+tpr0Lejeyt0mpiwWblJ2m62GOw6XVQNvuBwM
T2sGJVkUkwAom33WS9sVUI5G7VLnWr8GsMtnuoqibLcgC1a4DcDvUG9uQWj0ImfX5mbmG7jCll5u
TXqh4pdbIcytgS5Edec0xhBG9ds0xwdRcEfT/hcc9uDV1RwOn0tJdSfRw4/Pv+QXHQ60XsThEI9l
2wf5qzFKQtZq6mJUVoIQIIKDZ6c7eGXtLdtQmyTOckrFvlBdhBMvYn0p4Sma09cYnfEboMvFCI6a
pBjOZdPvMMXME7dnmkVH5d9x7ywWxAGxHW70eg99AOLieLLcgSSA8Kt03RFhH9bFp7zBXLN8e6F7
U7bf0B1G66ODvTdJXnOduEf9YJmk00jAlAqUjJCR3/IAeytZ0DYNRAQ4UrIPPs8G2EXJ8fqi4a8/
ntPbpnYsi3Gid2aWYjzgJevzxfUNF+75eUxesXYKYqo29776AWElEYiHzWwEGNGArXN7P9MAvCP4
sEYXDelSeuCK0NE6Kx/bglaMfhD6RkgjTBPgShjhwzg8E8GXuVPv83RK86DGfCg7fv+60Kb1M/ZU
dq7y/ZmukJ1V56T+pRlj8vj50J6Cu0LI4VjM86rJNJ3nsmfMVGp1SuAm981OHZFW5RfKTubSe/mT
PEGBDhAoyJNn5PHjm92feI+jZn2js5HYIXPmxmOpGaZUfOS0IaawEpOBKK4txK/j8Fq0AfMloefS
f6LDZHG8fIwPXzze2eIUMpnTmv7qcVJsx2RqoO7pBQxSnPvKYL/6yvEqwNblcd0uIXtOgmLFpttj
9+GSp1MpMulBFNpb1dWwNeN3RmbGKfoPjH1IRZEWCMYmS8PjPPmdC6MUlmmwwPzvBxzV4491TwoU
VeOAEYHcAvmqGO2mdDjXPAXsVEC7AvHavgsxjvv4n8TuzSYMVuuRfmt6DPWmxLp098H+YUjntPYS
7xRryURRKO9Zow6vbsMPmclJupFqRttsw1OEPXKEM9mRhEzpVMzslAIfHJ3HoNsyNkZGIpOzkobw
S/Jb7Gsg9Sy71JodtUQLb3Mm0L8k2tPfbYDWHVG/91pHWW+KXSq16BN1g7AUU1zsRCMjHteh62qX
Lo2v2iFZ7Y5j7nmknO5tbWTZkp/0zUUR3q96wD9ZhEuSuUfIC1lzt19yrlD9UQRG1wb1hhWClNKb
2RbNSvNAQ+36YxJ6YM+qh9z6m+PzYbZvhGhEHDI7XKhHOMIGJ20aDT68YKV0GjpmANR5aeqaVW7N
Orfg2YP6Rjt6pe83MZJGRsLVk/0j6VAf37iH6gWrU7VZgvNRkpJiv3b4bXiaPgwhYXbCX8ZYqnuA
MmoGrOWOy/KDu6sgan643tZbu1g9qiC/DLDbasWtB0z0kvW0+LHSyd2nthIwkIzlIpinBTCuTMoL
Sy4lizLpZhS3eYjdsmljgHlt+cd+/uAl64+cTKLrSyAFyqC4bgVGVTSUHLYXO4qezjDcP/ob5LY6
e1mqSX0L+YX3pYOBFg+M8Hcyx+IbLdDn7PZR7SkEFVlUKTXKPAbrrmu8hUtzDI2BjbIKAOwCC0c4
7nCZxRBKILQg8JhgsLF27RKVYxxZhc3QtCBJGMLBLIryffygtvLXFEclgoN2Eamm64hYdrN7nK7X
78CQWPQy8/LOMDYQLZ8dZw7qNKrw/1iRVqjwr7Q2JCK/lKBgvK37jTL2jG0WQCoB69UITi1BDH/n
3CHAD86g9DYQzO4YfxdmSFMOxOhDC4cRauTecCZ7Z1r31JbLGuQcilz8Zo0JwCByigE2iiB/TPb0
GX6UNmDkChldWZSSXJhLgbR4l5Ft1pxFbSR33W5/3Vw2z4DCQJVwtfFTEF8YCZngkuG6x1jpmS/L
KxaDrjIKo2DBPLcN74wcrd9NnxBDdNhyIe2QG5agwah5kKH6vOhmWsuqRqj++7YobUNQgHTKQsni
W4gsF1C0MC2a9lok2xOsB1UcNkjNdenxedO5B8rVBO5zEBa+E+JF9tg2ZmzOTDSiSxLIUJDhQP9B
Eju8TPP/pDwBkAz6TZJbl1kmlu9yfV7Qbf3SDCFp6FyvtFBVqvQZoDD+gHMF1uBTGyJxqwLb6Zsx
wQaNtqVaEW32yDgW014mvZcWlcRV6RdNr/QJIosVWsgoGFQBCtS6/u9O3Hoxpey7pMn9AqN1lJZX
2mwRkaoeYPt1djJTrFIrMVLhgb0uoYftPsPpBp/IaysG7Gv4AQ0MZ30Gba0BE/AfIP/FI0G9La8S
Eum9yw1LhXFCf3G4W6o6V8aQLo+ZmWWsDTCxDdmSdBeNPAENjuBPaWadFFfOQBG3hZ3TLRVbcPmk
2SDXCI67yPuVUsJaK6JFxaM87+gutc/2orMWJlubDcQ3zG2UF+wkO/DRQLjN9ZrXwz5LiIkCjbH0
UPhsRO73Xjq8here9U3X8iBjl2PhI5SgdmMjn5mObVAIjJ4xO3xy8FNQmgoY3A49VRjsWM8DSBWW
TI3T73BqSPfJOBsxRT3wWnJntYpL4F5yjs25ILbeI1acUuf3ztiOBf4ULLJEuA7ELvXBr2x9s0m8
47vXts0AM2hKCITOc0zY7APltYRxjFKYAOIWtwxAyRNHYhnDJWKS68REemNIMM4haHC1Gom9S4Ay
QfE1dN+810FUjBDj2iHnKTAZD+7qRX/EcfW2S2LQv0MikfWLHrR2q7P4pRR0ba+TECO0ePU10P3Z
YBGv83NeVkP3AKCQ1aEizTFoqDmVvs1+hMuyvoV7uDH4pJkqIT60dAYrIr3l1s89jBSliPhjA9Sa
gTCpToH1px+p2v5sAHW06vzO0bxoCijryCdaB3J9EjeHqawHZoCVgPREEAWuF98DfCi1V+ZbROw1
oZxpciFUEaoI3uTGLLY2Q+mQNPD2d8b3DZI7We8E3DaAbAkiUByYqD+KXLaO6468qF5JIQZFx5gs
EZ326N9Ih5Twtg0NYhhh6+nLbFP89qWNQffQm+/mqJFCIlGqcXDn1e0ttPpUvdK6twkpJcfXYRYX
APUd6pgXLAt9wtwNo+XcERn4TLhwzsyaSXNKdjJX+2DmyznLhLSuqGbC6L6LcP2HxOZo0QjJfKvu
nF9jDdEbuTbbVCrY91vBTNBLjfTH/cs34Fy7ueQ04s0Tbhp+t+lIRF/liQnFalDPOMKyIFxipAak
Mq570dOKudcJlXBhqpqvO/iwBgn2L+DNFUGGgpNsD8Isq6JtR0e9lEmElZdh5Xu1xpCxPHCaQFdm
e/reMu+tuioCLvGb5kW1/7Ipgoa5/8Vuy0r6Otsj+O0bh1BCjUG3oc1SPTnVUUmqYizZDjG56irf
B4s3oe4UBMfm+dlO9OuOProo4OK5IbW1QLWG5QFs2HVjSQUJ1FhnhazIQJVP8beM3V395mM/Dvc8
tEcbyG1pualYhuRfGVLlrZSHcse3t3TPL8/f1SkL1NUyAH2jGaNzdXyK0k78ZBnntaV4TukR8xVc
oEAx/ErDokqXo6D7ztDAQsw/KbYWyY3e385vbBUXcc+M6rAbAHlWwNOuPbTkIRyVcvHMYZ4ksM0t
y89GT5J9B3Nyv9YFD8hlKP8ASKvheGZyHy6j/4MEh61X33bCMFMaz5uC0uAAx+I6h7vX/XJqKNOX
hVF2C9A1yzEzWhFGjlOrj9yWmHg8MfNMHxQu5P7NoAMlPmelpfqxZJqcqgQxpZ5NFAJXvcZeQMC7
JDFQI7kCUWi2lwvmCGyyNSpAXrUaNyadBNQt0lhzRU4xXV4zlgkJjgqrKxxbETFGuk5/uxxDG07x
M6U4gXNshy/BhCSpgdoxRQ/3XlN4YvYD4Saqn3gBA5raNSxX6x4FBXl8z1rt4lcGhO8BMTaKj64M
NBZhPkjesP350v/qknBdFoLcVj980WqaVjm4cuYT1o63JhQXEha5m6Z84KL5ouNVscZlJ7IWSZSb
dbAXOOc2Z/2yhmJOpyT4Dvj7LVScI1YV60R2NdmOi7kX2ZC+8ZjyVHm1ioSD8iG3SK3raJf4+aZS
m9wpLbL/XG2PdTRJxG0dyhHXPxn+45Z2VXd/y5tVRhfEV8v3cPlmlgLXsQ1oCidNO2pYyN9RJbuT
7yL2kDIigv4VXIZD2O94Q0UXg1sMB4qktRywGO6e7p5vgLUi36RHyTbRC9LGYVpqZS2uXuISGzLD
0Voc0LHq3h5TFM69AAUJp87GlPicy2Ed8XTZ52VuG7k+h1p+OcmX1mUab+Qp4bXPeDSQ36dvZIAC
kmx74ZPnYfsMfDR1tH7gc4N6SA4HOox4CfS+8Qyns+j3qTp4YTVcxrn+BfQd7BU9gwXMJW9XHTu5
SNADbx8DqMADBF0vIDJsiQD8qm48UgcHQbcLhjdENrOZTlYLmO5uyrlGn8lpBvOgpEMRGYwhjb1N
zeyI76Y6JHcGc10ntIkIbkPF6BbVJcYQYoTos+PTu5Jxc0oZ0nNMS0PCzIyAaCsCuVStC0K7TOFd
1tFOgFFQMivaiXt8WcPWGSGzPXNoKTgHEbWJLnlLMKvF2vAHdWfTNaY40ZkW//vmGEy5Bybi0QQx
YZT62Ljg1VplMpVobQ3sQIYmrQMY0mVhgK9SbiiLx0fTexv72f4TmMjHvbWYlxOP5VWcjs276p1m
oa57HNw4pxlqxfWy4OQ78NUHvPpqE75ah6jQGX/yJ6NN9koC8D+190mwFgX9exxgbGN8YJp1svVP
Ikgh+MBChJz5qOTm3vRaQW+LNB+Vel59vzfNqlMKQmbmCUAS7qH7Y/M6OvlyBcxppDPUaq9216fL
Z8YjYj6+iKu0l/vJ1o5qex9rNl7YzEZIT2DOgjUaz/Os/3bw66xgcYLl+reOgM8EQAIPrKj1hr5M
QUVp/qTd2yxDhH3Eu7AsTPGrb3D5HXD+AzR5CyWEF/ACkbz79oiZaATAmKa2SWVJuZKfSED0LLQ1
xVo5rHLEUATlzJYTZJ7htzl8JF9Wtr8G5t6jGFy2tNIZ4jtYP0K2Sv6eNa4oIZmXZrGlWafDpOkU
Eq8bqoTlnWUi2/saSZ9UInxsG+mN91/cLQMvuxmiwKSxgY9Q5Gc8iJAES6YHEiZuIHAaG0SfLtKt
ht/8NU3YOcnnYpwV21E1N8aMdr0jA5HmRbuuRRw2Z4C5YSvMlLCgAMfI1YOvrnSakP/VvI3xaVyt
kD7N4AiHK7YP6kxRF8rUWaPTGRKDzCU8WmP2gbdNAnn4ZLfRk5Q7QWvhj7r6HO7cb+MgcF1lLdLu
2yRmzxMLeXyK/4hhB2ECYOEKxJ/Y2F8AgwujBJMNTVz3OtcXh8jr87TiJshXR/Jfc1nmi8rlQEg4
+vHPB0VScjP3rlk2kPm1ate4TzCsYt1zoTafwnqlAPyr1WfbCqr1Wh3UtrgD/JcA4CKUI4n8C8d2
AaPlgaUr/reMCQVjAHhrfTcmFM2UFOoKRglrtvDhNPzy8wrKAFYRo2C6thv0o549uIfzXNgdXaF1
4XXUPwX/XuqVGJbHprlmB/AobGnMZer5BSZMIWq6+93ZkloqAY3yW1tF6hAG41t1wsaeD4pdLmmd
6cyq3NAkNysgUWNekABlqA+1glxuInp4fn2JdaM2iDOru92RcRBPoorhJKNZAeM4OlHaowRQ1bqo
63GdDWLIoevoy+IjqJruwreiMkUWnbnsiZ5r7pNYKX5awkjnMd9aqd+gyIedvX7A3pi8xpExqJrw
Qyj3NStRq2Ui1SzetMFCkATgc0lvJ7lH/b+adGfe4NUHGLQtJG9H2R0Q3Vx4dWrFEf0aH0ZSLmK0
P0RppJmvTBLDLXeLo00MXsPokMlczh+2KX+KETPfKVw2ziyWjtSpVnGTTdseB5vM/Ct382Umff/R
k47ojB093ZhY3GVUboNVt3Wdyw/pRW9SkyaIVlH2ywSfdRQoIHATX7JJDXDc0bk60VrrQH6+zZL2
hGza+m2PkPIc2TDnl9AQlLunBteSGxex32Oi81M24XD7Y25V2r1fixW9/FYZBlEDrvQE1Ebdli34
Ukgh8Dm7UjG/4QP1jcQXZQoOiAfRjJDRybvtFN3xTn1IvqvoTwyRhf0NvWSkpWDhZGDgM4E2ajqr
gZActFtOMO3tGeHFGEesVV8R4/kyipCctL8E6vxByoK2LXKrQi20AvMN2EAUcAyeW4BoLEAoEjHx
qWh80XbPL91eTb+UFDAZXKVI8RiJneL1P+tWZU5rAR08xqqF07sTSUqI9pnyi42ZtDrQzJsRuo0a
g/M1dNa1yoc/jrXUj9TYaWdNBkT2F8Gsh0Q91nYrnk0P6AwmOVU5tqM2oaU2ymYlWI5583RlsmTn
qsWJjWtByW4I/y91mFTC238LtXstoUxjpAj7Zg6dmedWMgcYmaNMDNrOpzqaT3+QcoixQ4K4OIym
Nn4CxV08+SzERrMvYO+7fLfee9yhXiSjIpVUkUlUfjjzx/Rjed08lint3YoZneS7C+UdT7MDzCNZ
DQsXV2czg08SyzBDr15gjwYC1xqu6TMaNO+M4Dp0kAGc6nLaxBR55Yo9yR9XrxXwNeMTYUJDNrKs
QC+QP+1aQoEjARc82lowHy8q2swfwaDXQglLC7Ra5KXZHInhmH5sCjqj7xNHVnX3sxlvJ7vbeINR
jzlgkbB7iRfUv28tK79NKWcA1kZtLi9C6pqh9ohNhBFuz3Mib1/RtC+o6u5z2SA5pMHK8/VZJdJm
4pDTDDGJh6AIu9IJ/iNPoOszc1MuHOmVMiZJK91bfjkFbXagDjZFuyaaxlFNXB/z9obgGnJlCjlB
IzeeVKNOnMr2ZA723XOirtRjRXEQIDgXN5IAEJLQwHzoDsDyei3swCadw0QEGd1SHBNmo/OJsTcN
q7Upkhdf7yNpV6yfdaVKKiRILX1NGeA0ScLeECg5mpi2owdcpmhcLBd+KFRTDnUe1Kb5duzOttpw
c3CwxTH60juXY7P3GB+P6EMCugMJg+oXEKr8ZiNMtwDJkskFaF1p1XYkNLllX84OLoCSb4cKM+gt
O2IOsJEqfghPDEWSGYoRDN0+xNut80nCg6IpwW4MQngFBMf4ha9d7wWZu6UYKQwl9q3MlY8eeA9H
7KHSSxLiexeafaF02AG6xj45xlOAGJmUqQm1CRll5j6Js91UjXMrSeZnRwb2ibxdiVmLHe02/GYp
+OWOV6yd8kbWpjxnSwrUKVFTBQlw9LN3xS8ch/9zzwnwgG6FX4Z5UPaOVEH3E8ZgdyT03Y+kMYzB
BmOQEwZsDPD5jaXbXEBAX78qOxSizWOcHhUUt7wM+wwheqIPpq1tKuFjjsug/VLKXpQZTabc3QoW
lGavZmUrCLcub4oDRCIBHZd4Twn9Zmp0o0kCFUTuyvA7wCk7fpnNySDmPjfudtBBlTmiA3m4a2Gc
wdWXtPBfCAGFsepAuY7Jesi2GG6KqaECx5/hlX+22h099ESWAUANLBbG5eqSgxmPhhi2ifgMYoAf
1J93vxVLOX4cWrI/chkazaBW9035sbqOjjY9zL1aDPkBuJmBGallnNhaXo04sH7Aan2MyI+DAD7F
nyEtz50qqFarlmx647Eym3+KU69V7vgtbR5Tne0fj60d6UI1X4R0WsHXHBU85mVHDdvtbW5SwemB
gR3VgSAY2tKjCaqoYiMRDSI8k6X7s4UJWeaoA3uq7PToM2RaKPXTurnVZbVjHtb7D+CEvx0CV2DO
EjunUgF4c6xtdZ0frkm0wkZi5LdVZQdtr62Z3Z8qeSfzo33sGHHa+LKdC09bkz9Sebm6ULqeVMRQ
4z3JHwMRpSsxOthMeZg8m/3HZn5QO32MFPSz+whRG5O6fs01qX3Yxs8WhC5MgyFtyZqzcB1JghT/
0iEP3EIkRgyl4qubL6CLHe44Yo3qraWLmUtVGyyhww4qBl4ZOXGuhTDxv0r9vPMqzvPCV0LIHBdv
vfmmYDNvPREVtT35+WAiKNS5TOmF8j0PIBcht2VmLW3xzlYxQv22cfqNY51hI0wphCTrSD4LPRVK
GcOxZ3Ea0uO4NniiE0in0vF96zDHwaZfAxtoQdIgBX/r6JVciqrI3VT7QNf39lg6qptvdh8qleza
nzHXn149q+o1RmUDw8TDndzhvjrrjlkLmxrnzmbiH0LWzZt/Xguoo2i34ysSHualjon/8XbLIjr4
eS//wt8btHt/8cTBmllsbAfxKrIpiKo4yQZ9yPAmHu/lE5b2gebXnYNzJ51iOm8jPa3GeALABcqR
tuo2WAZbgdLiaHXdPs2YfyOMb9KGbIHESy+44Bw4KWnB3sIIE6q+7QtWy2dYMuuMdBM+Me+6rVfK
BpOfrt2oZ1vqFkDF+IRH6TeikNUmMW3uctG16PuFFAu7uYyaBWptvdQoU+barY68x6ej6fxNrUG/
TtPO33Qk4d0DQMACX5jSUoAtSwJm7i4zZzsJ7ERLtQRwfvywOXZdo+S5Q5m8JdXJVtWrxjSh6ogc
ieUjgTo05RAzZEbIQuqU/ZN3KY5BQ3SAzK4s01/Cvso7Fa+WRaw4FHeCE5fhV1zM7AVQAha2B+rt
HIpsgsk1gzSJ2fKDnPHCVqizKZFc/hHCPliz+Vh2KopHRyN+Zl1EyamiOfNqG5aT5oBrBCVF9qgb
KbXxLEMlOWPh2EzTy6xJ4jiL/n1C+35/MrcAoYMmHZ4fGgXnQNPsfZQrQIEC4gHDtqOo6FdtCCAc
3aXNOm9jnbF+dmxIJ8FPFW+hIjnsko724nyt6QOGk9D2xCl8k30xpnpUsCrRjcWwILSmcPH8pzA4
iJujZgnA3Jfz5jfQbXRr6Vb49yM8DdgMMbvv9dtT6U18UV/bLMYX5tKrWdo+psaQJj4G6ujgdpBT
/3V8ghnmaedwumH7XppBANwLMPs0rF/VOL9PTzrB4P65Ds8NUmOjmgjoJEq352hkUM8gpC7zeUE7
4sXbD12tQMpBGepOganN63JyPOAkKJHq4g97+JEyH9cAu87Iz9VwNKAnIbyvDbbQlRabpKes2/9i
Uy2/r4tQNYQBSADajMH2jU/P+1tjXhz63WoWVCvtBK9bl2qL0msUAcI0hgo8OYQx64yz5BkSKzc4
86/QtcnGZj0YngIY0QbR5rjRvlFsCyf919BBcBkQ8YLz+nNhu8AoSqH3tR0WbCYOBIR2DIGJWxVQ
GpJ0Cn3pugXdKfcNzPvGs2cceHvEsQ+NaRaYy5WEymDgGmSEwBR4IiO7Mhb9bwcqClIz7wShxD1G
GKCW2MdgpOEWXCBquaPnjJJrbjppcuEgC7hxkwZmV2+j+TwOrsjWdHs5uk+MbC/vSurqp+P5ZQor
4g+VU1yvVIegBhahTcjv+zLKzP8yGqd6V6mSfxRVuD9tXFaZHLWt28mesbQ+D0s3pKDLIlPjwWhP
CFOp3WnmrcQDmWn1HRAOTrzGSw/oYA0I3WO321PVzN7uihwHAWGXEktUTFZAx+E3jA36d9yNE7RL
BnVHX6ECizxkBpVho5OMOgDJeSagq+V3t5ZDy79rHBpq20clOPficFlGmsiwHmbo8jw/xFG4pZbb
z64k6r1NvHXexKLvfXz+Ogl9FJHqon1K2DS2/8DPAGEj2MSwgPbTQIZVN8mM4cmJifjRnKwE3XD7
mefs32hCGQRYepknk773m/ljuaL2vA2385sXUtJfaqtl7lCaPZNIs5A/Kyeka0LeMGeVLKFVCfTY
BfuqGdl9HQdF+993NgiIh0yr+Z26/TJv3X3gkatNa0hhY6oIiDg74oo8yxIqNIZHwqxxkvpkbQg1
r+Itfl9nlp9sQZbvXtGYle5A8bOviV2FMxFbIdsw/8y9jdfKXT7R8EGl4N6s+vulNIfPw2mP4exr
0WALBkvSAFHv0q2I/1XV6DW5b/zf+OfXTjvj8TJS2r7/VcGfXhL6VvqPVYcCRr+Pz6tq+h4m1vEX
nCHG5YhTh2CtYv8MZW+NtF2gGV/9sj+g9IBQDh7JdRxzwk9U/Qv8+9ic1hTg6KPA0yhIK8NabDY/
Xf/lXkletnIhc+w7JVjCATLsK+sZuM7hxYDyAuH67EHY1sQDy1/E5UKvsvNkPO1SJQP7HrCFg9Nl
z9JH36LX80tujaZQs+Vx3m9lmLgZi05GD0okyVrdg7BKUbLE5VRhM6V5SKhYhJfU3lyeHHix2aFZ
8W1Tzepf5fCagMf5I0QH0sFfDKP0tvaNDoyY935rqGlevmU8FgV61cNmVA+GQqDSMbGCbjoXD2jQ
0vAOwUQVv8INfCBt9ptrbJCVpHY62Qt4ioeM7i5kDugQqUqJ4dbKVkim0P9LSDwayIY+e9w3DsfW
SnNM31WjYWa0NySpIuwHC5Kq3/oj+BSCjQdYGJiZimD14JB4wAkv/LxiRbp3bbh1bJGmLOofp4np
ipKQ9/ku7r+nL8grhWK3BGkfPQkPSuk+SEsIpm1thKbTr5vKXaewpnyk18tbBT68imRnrkgHqKZp
WIUXc91Zet6B1Kshu1D05Zst/fAImNXNeNq3hgq8G2zT3VwiO5hqMSDmgi5UeV77CK1n4l0huF9Q
4LaTkyqUYv2kcRjMvfRNq9xeOewrTJYH3GtyW7nyTlzCkma/v+6PVW/8yUXUWhZutDcsHrGoYbCY
pL18o0uEKppvatIIwuQsd6zCFEeOW5VAZCsdOscxynTm0UJmFVKsPSNsZgKpEXi4/7yXnTx+gOem
1eHzhpHe6Nci/D/BOOuAGtD2y/BX3HrW4qDHYGdW6Ag2KrKfb8LMYTBSqsbzZCUYDEzJv3j2c3zj
vNh/GBQNslyZgoXe5657ubyWJ47r+qWUF07hjB2MhNYYts17E259+7UfxPhg0g4qnJRdi3waPEbX
70pHeC+KCeNaWMkmIJN2GuOaT3Yo6sJoVZWIH0mO+6UzckeODR7KbhGU9y+FOJlZ1Ig2gl7lxwLt
i3FcgFvoAXr8Ogazu5DbLHm/NIvDzSTRJg3/+tcBgT3m45p5TLPXut8PLLoQIWVBG2Borr38P9d+
fTeu+a6h8QDNugaR3hfeZCAbM/9QaEnbOwms3Jlpaynmvqa2ny+5iS0oQzNoi4WVf18QyQQRTgBZ
H3xiG49PDqqpHU76mKlnkhQwkeCNR91EFIBn2Cu/ccNozCIK+kt8XLq2qHkn2ievfvylBnrAzc/6
XgIi8scj05kKte2spo9z3AKFMK6C+BUHUZ7zymmW0R2AGU3ju3zCi5GJ1ItIA7br9sQbdisd+zua
7g19/KWY+I14RydvmVxaiopFUzgT8KUyPJ0xTIEnLqoM+QySlheYHIgsoDdVjY2jkWt5r9tVqWNI
sVQpeB6yH1Nrz3jY4wPt6eTW39xmq0v9bHPKbRMJu6ACC9b0KbDJ5EYUtoCt7i2yeIsNvHczoPj9
f7kmlrl+/0USquFrw6tMDnryqbWIP3W3Sd2Gd5zmTZW47F3Mtk3klVZ+gUKiHB63CpjO8qDcEHDy
GbLWGJA/v+wSW/oKb6uz71c5a4auXEJdZbXf7RyYf5+vpESm7tsnCX2BsCgTdNLb88k4Gte+v+Zo
T0rwwCVX6cEy6EFMt6PfyNosKfzwkGX25qdiVgXrnuk02vbm29D2lSNph6iIXMCailAMdJAf5AWc
Pngs4ffuOzrn54bulDmjTmWr7L/2mShK6dlw/RpG+MGW2zrOY9ttJDw1m6WTar6Br613lQSX9cgC
4/80hPjUJJNWl92L+b6e4QRXzF0D8WlT5mFmI/sGSXZuwWyZpz8kU11CoYOEbg51DV5tTMCtog1+
Wh2OXy0XdYYDaGuCpwyq0l4frAN37dJZ++rdNbsBgsd6Iw03NNbAL1YPJLAwlUo9/ZXdhqGX6cS2
2/UG5A/cIB1uzkwf3Wzd4G38tJsAgwVHI07Z3mEebOUiGtJ2WUjntm75YNBlwX323bGkqKwZ6uhc
U/q2bxmC0vEn21wRa3PrRD2JJmzYclGPd3VmBW9/tnPiS/3JobgUVsvaIySzL84maaYk55DxtbSw
aWX1C7WWQj/PDT5meqr03wEyYPBKWC8YDsWxCgDNTz+GYVBtZ1Ae5d9ZCitEO8NZaEnwDU5yqLWZ
6XIiMK6kxks8qmhyQOK5XaoTV81Wgux3XOA0GlVNpAPPs9Uo9xPzJFMyrs/BzGZPiM/GPK2vUVST
slWHXYNNcoC3fwS56pHZxW5eZC0OpvWOqXpXASlrvAXDLOBqEdnD5lVFuswq+cvHCVN49bDedZlZ
khym0F1cgjtDKvpjbD2Y+wUBSnfq9f3jPYyteTr+lHDoOIEugzDZyC8iBBRl+6rBPpmYAi2/lfEk
YvCvGh2F7/k8gB6/zd3U+8pbiqYkEIU38d+YHQLYy8eQc/ZNnNrrRoxLMxhyfXYHmiJlrSviNrGb
bRF2WEymthuvIMiTwbCIw+zO3wfVCsyc7IdNIFjZ9IvDHUfMsChGvZl/npx1ZNL53PzzdKTtTPcW
TiJsqcisZWY5CGCku1hPK5UFKi0sy204SFrt55Evtv0VxyAjNYG6LooT66gX/kga+8bZaYjUOT2k
fynr3H/tggDTI6wfURDGMkQph7LCrFMpTVovGEn1/DWzQQd5p9b78n5maBfl+/NgzVKrSJM1/60/
vln31yMIUyvLnLDbfqddwv4PD9fRRCvlsUHbCst+8GlEBxOSPF3Zj+k8QYP0osf+mt0qvegwwrOd
qzqzBTJgE1tYEFJ4ePpadv2yoqePLph7BRv/yM+dT7K1qTiEeqQ6ZqzaULy8pJFftWN1JSIoh6/Y
yjFiEZ8fzfsNepRVGT4jtAdW7RxwIrOuUrxGRUWRf2Mb0MvzNKJMq7fVchHz/gC2ISZaAvHHum6S
NgXpWpGeuJ2J/M17XSp5Mze8MFzBzv3LdJ5EtaEdffRgvy3wXxk/8z/1YlIUecPVCXb0EjIneACt
H0Crpyy3JpnTLIAiIVTu6gp5sHYXYwNosHzyGB8qC/GCVmP0OZRiDzwQAveE38+awGGJwBnGNnjx
0Dz2ZjRWnd/I68OLc8Jg0vI74tJNb8O/zj3BRcGk3zZZ7O7opSwaorMfU0VqT/D/XnzPkHtT5UpK
YTu9ylXxIHzrnqX6SmxbnNG1cjyh9fBgFXnJWfZtxjm30zBeWTAOs56ysLVvYsFbZCw96lES/eqx
roRvwFtvHn98X44i2n3Ug9kowYcnbrPZ1L6P25HCKETIQZ2aZiZ0qvlOIEqXA2KF0hZsIGVQa696
zkvRJr0C00/kmoDh2s3aHB3ULrG2mj8pkpzKi1ERnalIKDiuiinGXK0jWuzUw2Z4GbrOUqZ98Cbo
lC2oHLMT+LL+u+KJfzgkz3bWfaiOM/BcZFUAFrOVDl3m28yoSee5k4W7wztMuRAhZsKeBzolEf3x
osUAXtbDiQexemb9HtPYI1YlDq8DoFgCopBrjPpixFdapXtKplxCatNqKWkDL/s9yKKFeOqWzloD
X3sf4d8X40HbX4OJa7c95S86FFRwlRrVDlV06QdPM1b9fVpE8RnnTAVtCSXDrY+z+zG1y95li8yj
lVO8bh7D46C5ilaNvOQ45sbpojUZ5nsBOZGmrhWGh53+DXT/1tO3S2sXqhNHDiNLdur3bdJHgbfA
nX5iPo0kjdcEA6W1OAhOjCnlHNNq1JBfJSDct9TEN7NQxUvMrfrFuEqrL94/9jXQ84i9V0xKNYJA
Si/U4wnwSsk84Cy9gJ/cyVQm4+XoS1/UXqM6CsdIA8hani0z/ESLPg4tRiNn1Mc8ii5afYgV8nXb
mCZnE278FqZOtbMG8GK1elHeBResvWl658p1eHAc8O4hykhpwA7uWY8hsZeEZ3WkjM+ow7Xpsnag
ksEudXgKv26i3opEhKKsu63X61i7Apr4aLZ2/aDzVsB9/kwHsuvGPmiu5YIwLbJlTvTZcJEmDnIM
aXDBM1T+vNECi8ERNodYfUk+PvO6yiH8gpNagkO0YCR94PV8tphbCtUZQtNaxsmku/tQ0R2LzHPs
tkncof3Kl6qh/Pi8A5wPJ/M0zQVvNkLu8IcsG/xAsJjNLtA0lYfGRwbMQjmviTMim+aT0hlJSmke
ziZNTBtNRfJErtzMkcom1jWeHc9b2JMuZJJAnH+2FlZS/1YtTjwUIMrBJGheG+7d63jUjQl1HhRC
Jt2j73bFEe6eyDinQ+AcgG8IyAFBWZMXqars4RDR3bn7ACMmrua8Duak3Y4DoRXdBibc1YCQo2gR
eKNHUtIWjHV+3I98TLY5r6ihZBSa3psVwOXYcWMo7jsZZHKV/w1aQ80QCiNARqud7YqpgHtbIia6
GaUIVtUoyW+uzJhAIwskpzCy2FH0BfFmQHBi4zJQepVJ4g7YuSqCujajGUEGkLUFISF7AcqzxTh6
LrBCj2ehNKpjOGdyMhioebJ9fr1IaXJFqZhVkHtca5cDqkE+zNz9xCuU3vfnXILepwXXmfb52wSA
ldVVYnTVA/cnvn+QQ6bJw/AoWtKyaSgZg7bKzpUEQK0mTfCMdxwgYBidu3jsNdW6szcrFjQFpiyf
VILrBbFhe4a2jo7IH85936aEZ5USPPOnhOj3syEqZPSlvb1rCCCQiNOMrjQLJph5/hXGpfg0UqJs
iF9gHRV0KuOeGStyG8T7fnY1f8vCbYgwBF5hZ/uqR1B//0pnlx8K+0e3MuYoOh3a/6AlEJIGzSy4
e6VMZQCdq4Hfzv0Fs7IxyyCcnr6ttmCcoJTCj4jIWzuZMwNWL/wYq1BkyBkSNuKrMjKeDedKi5Nx
6DJ3GpMl/NuYfZG16zWAXC5zj67np5pN7hlmZiqWQzGhDx46KjEqWsAIZIJkbUqJv+PUjOLfuZqE
5N2LlIrvJvflnapBW5XzBSL24rs2VNER8IMNStRtdWLnwXjA7jHaJiDSesMzniYr5DEHukVBax6H
rWhvobixA6SAHK0zbchwlcHegtSkAQVXcJ6Vj+suFJOQHniPR3CwxdrSzS/3/W4mRonldQYz0kVQ
9lVFSQm0HN2+NXpZbI+YIW3cyMgoW77RdzpNsWUz+2dGWXC4LL5nCnzC/SEIx5ZrSyF7aIzS4Yvc
8A18vGalo07wC57n55DePn86poJdiFjJe1q7kAt3vZ568pppkCsbVKzD+X2Z5BpFdjLTyLNpRnTp
oyxX5ddIRX0Gv125mqavQj2Vnz4CLa2eLxt/YY6rBvFJxlI6ArtIwCEsR4pOYoUS3EbjARG4B/+m
iDG3l2OjINGqgcXTUwJDFI00WNFPVqfGDm0irgUINfvwTmbBIsXTPubVFRNa+bJ2zJ7lG+V8P55g
oiEt/M2tM+VEa36tV/fC6yS7Beul6k1C/S0QGsTMXHutKzuH+H5RCsalkUm/PTAnXruVDP6hyrQg
yalFYXHtfJJvnMLeBoXAPGXo3DVSPyyzUwrbKSTArOy1TpBevs0B4nb+5fOsBEPRqYYMXbiGWn7E
9Ps24OSPJMobg0dRRWRr9j9vuDMdIYEcpXiHGUYns6dXyxDLDhfsqe5WNRrYRZkN7szZeY5VGPU8
ihpV8kob4BfwhNNHPEfl4mcQDKNOEMPCsbG3cFhrJ9gVaT/mwYmsrF3zDILwdBb6xtKP2cNjn8Kr
YCJpVEjNhyQzP9WjqvSnE26hrEeySWvLMe0p3424WFUbqEbmoE3DFcyYoKNYLG6zt5xJ1SsTgipy
bvI6Lsyu6wGVLl2tssxemYB8c6dvoWgj7jKpw1W4hl1PhSWzPHs4oNUaZzVDH3TEXsBMucWDwOEN
nCAfLH+QXICCkCXb/nEn2TTf3i44PDmFlIbQ75Gskt+7lNjceyfoOEj9m0WvBXEO+HAOZmx76fVM
UB4L51UqgDe4G9pN/s3pfrFShNtk2Cq0JSM1gms7OCdMRFlLnNQCXdUz3I0YB8gefzYYBgViLgBY
t25ZSGulVNbsHrTRPin1b7FzVAGb2JPdwsUwgFKhxZtphO0ocOdHWnkVcDUwV/Ff4Clc/8WmR5h5
udGMT/QiU7uLtcp/wkugkdSX4lXYFyD3wbRDqSWS1hYQkAFhQ28+jt+z66Qo5UzgYmawYhPVSJTK
Emxu0wkh8Udw40lth5gpBdGDxl6mpTKQDhV8XnDW7QfbRRN6rLyx/PS1zNQqAU9Xok9XfzYRPjya
4p+A+7nDyu6Ehtq7/ouzZ4ySz71v0ybjg8x2X2oPdzbBjbXxs/NjXxq97REBajN///AWq1BoWJ3U
iCtxwUkuR7VEEhteWaHfQ29khBOjfaFjL4iML1T0aoy+RKplZ2w3v7TAXq6oeKAYLC6tmZ5j+QWk
z2Hon42XgG4W1yUedasfMxnGdPOTpLE8V0KJIO/MqaBS7ZpcSxeVzCB5d0GBvZZ8A0AE+Vg4QPRq
K0pR1QlBCPitpCYPGxc+8UuDB8+mUUjQ5M70j5PPcH/8O1ynAEJ/FGhBWBs2NELBaXjg6Umf5U/d
p+3dK+KV29W8beXGB18UgWq63+HBVjf9EX6ofdLONTrjQEEN5nSN81xhZM58W/5kKlvBH2AaVj4k
x92C9MBdPgRHCYKIcOZb+alryVdE2rAtN1FhfNB9954PB4UwJ1tFzzzHQvn0Z1DNq7d3WtIJPr83
/7sKqQzk4Mowe7hOj7nw39gmBt/N3AAsEr9Uj87cHFTk17l6v4DleP0v1y5kWp9mI9OIrC1mkxDm
UTE8DVNc/MSSu/oNLKrv6UMG2ahRW7hs9Z7KwywD2ZaQ6rm0giVGfUd7PYefQVvWM7i0tKlxSUe1
DnEhfpkPkxLrh2kmTsU7avf4QAiNOOZlTgZx1Bs8/+sp9/jyDRKnoI2jepKSk9G3V8++a1Naob9J
eMjIyewgp6bgJh5h9YWERDDg/F+bRoQxE4JmNawh5y5hrDAxDmp6VZguel8L4YZWwLFFrt/hIzQd
Z2vskGjNBD+D4ID29/0eCBeWzIhAIQTkP2XvBGq84O46L6iWrpn7ICtSFYoFvrJq6ApeVoQvUMIE
7FPEHsy+qWCoNW7lVegiKFYqPeXUzqkOonyVTvoY9RqWEOZJQWD2Ha/oPwsz2QVHxkThTvY3GXgU
K1KiLfdxD+l1b7YE9tK2WfQGLKZXbCcawKF9oK+CSCX1Q2jUS5W2WFJQCW0fGn81A0YMUNM3B+lw
GCK8jmiwExTY1LR8+SW1pEKSxCahMNvFpZAlRuQzlSGS6KA5yrAtKxXocJ/yQCP1N60M1BuRYdXM
u7N/OeVnE4jOtjsfGQfmwpl2LoQODPsv/1ocM4oVhD+KbUSEEhxn/jIu/4xDzJjgGUtabjp9JUVL
CVFev6dOJREsjIMmf8xtXB57Hdpgm0BT3eQ7y78SbxRLcsCLf1qzHYlJRha1lKF0Ktsbq5QjUyBl
fUN8dKLJF5E3mndEtlb3Ite81lsEf0l0hZFmzVM0HSJyA9tlKnlQ4Q2K5efH618g5Lh9z9j25QnY
P+iKGEYkLxXOU/11/vjJ8iQnSA8sInI639460APNms6J+B7KPXAbaEuha4XkLsv+cFcc9p6agDyC
qdMpwoxdmFOX7cmvY7Whvx3ht4155Y0gMNNa4M05Ppd7ccGVy+Ix3hWL+67RKATylNq1hVKHpFmC
k+RsZViRiveVam/J2xbTddxjaKNuJX4hMMQaM+OIZMt8jLYK/iNgvDNpOzf0ZxTbB7UMK/i3sd+B
lOG4tNs9OkgEtj/SPFD3iO49fJQRq37WLvJH327LwzhVb7PxGXrJKG7F662sUp/vnpwaW5D+xKK+
Rx715eeolVAMKUZnZLJRY1r4Trm/aVGJe5nAJfzNQhsNk9q33Qcc8isgmQrGKGEVBRexEWXu6FVL
5AyjiCUEH1CCx3ej6qOMiKrCjjNUfcGWOkoX1bFpRDVTEL5Mqlix1cGj+JEScRqg/u/qSfdRbjMC
7UXOGpdIcXJIWvQp8NAPsFZpq97gQnYjrRw4AD0xCXjTI79oQaO3XZLB0EmWuVA9D1v+fFSOs9jw
hh8oCG1UW8/02BqBDfVN0AVECzfLkaWl6Au0b1tKQ1kI5fWB4fc+UvfsZCGMY6TyfSC/RP9DklWm
Cbk5t9FuZglBYLsqooVJF087KN5MWfJs4usGDtU4Uasdt3tyH9fOghMeT4VgvCXfmjw1nP4xiIuX
cFsquqeuvV36kiVkgegnhusf1NLWfhIbQ972qZOydWpvS7C7hAIePC/5W3H84Z4+ltDH+Pws6cp0
bGnO7JEkHEcBaVcr82aE7LhfnCORG6InTJfQPIzavRKfDPew9CW4EPSb1RLG1gMEh7BROAjlxt1f
mIZDpVFmVIETRS/eng1InlPkBV+0MkPrCBT4TkO6PKbxw0KsWYTvTipu8CMvgFSotCwCHUAZ7Coa
gr9egIG02ERoWo87ovTRj8OzeFXHCv2NcZ+PkFbl24Yxzq1t5onjf4AQ2nTK50XlTOvtaWS7BeU6
j5UVXBejiSxhv/LqRPsmERgD9cfM7AUiYWXMhTQkzzcQaNXiQj3JtiyodbMxKzH9g+WcEdTnydbx
ISGqirFBJqQLLJfu/Weub1rzHzyfRIo2rVpdO9nA21kJO6tj43xbJkvcZXpfI4w2Ag4pOOYki9kh
hdJmlGxdy8E0ByWnCKG96viHs3clN7VC7Nhey13MCSGw/C7ZpHLyGyijw5km8aJ7ztpW0t6jeQ9N
IQhztLfitxDJwmJhc73/CitF5H8fk+ZAUZjEUQvvOgvpLpF7OJRzznvMiOfbfqCklO4mcsrLlizY
m05Z8mi0VrJ8tyMBLX4hNFZC7DXoNsvdfGZtnKqODmWnzj7dYKYJ+kOXVRZen5xGiPA9o8bM6brJ
oNUvc5QJm9E2RvALAil+0XX/CCZzbKPNkauYXymrKONf+Bk8XLE73xyzIYB8pO0bWaW1GKGB+AuM
t4UfUoo7/bfhxzS1nvSFxEX2n8lEbZuLDI2PY2wlY9JWUUwImiYhoWdUu+5w9voyvXXSJAEPJ+O5
OoryTsUZSf+Qw0q5pl/Npr7lqsIA0ru0BDCoLKoFM+htpnN+RfCh28OAjJH7TKrbf51GBRDPA5k1
4uNy9MY14aBKKXdvLGXSKhi5ufZvIdvIMk2gDCCHy697ABL9sT7RL4kEC0iPziKEeZCRIBqVMzqg
PxrF10Ok3XwAjO/A+VbWM7fsXQCpZPN30EjsyP3ebOekYaro5QvqE+1mF80vZWCLxsJW6QsNe30s
TYqvOTOy6bjw9XgtoASGrqKQcNbXafhEgzbwERraDcBXWBEkrRTwc7RMM9FLIhMMcQ96zF5neqpn
wGECf6SNM/Grpa7ntN6/p27SWPsupSZtHzwsee8U6kyzMlqkvYsSwtlPZ2ZYwruVcxd+e0gkR53k
4q8a9t+utGhGO2gqGLoz1CoGfZ5NlqD8OI1hQNGCTglglxg7oTUzVw4p5QHrmSeTvrLpfi5IV9NI
mGDbj/OtJE7TuLqgzKWbW9G/kjb8YLF+ByKCLVB28dFxQEBYk5RG0vP0IK4tAwOKGCdym25zNOd0
GDh2AWI8ZK3NsWnNFz9ZZMIfZ5rh5BF4TOCK/g9DemVAf6MqlrUWwdJdn/IMYjwwWuTFzQAGvCcC
qFD2l95P+BAs0FXtD7tI3ZfwTcliXwCRI7/cm9Sk+3erxFH0CNL52nhYgCsaV/0V5Z8nNGXOPIm3
D1nFbw/piqorze1lRty/f54vsk9wLfxLVW5bOlkSP/Ou2YNLfDiCeAhxJ4AcHZ/6zU1fiXVu0gRk
mdy6KjtceYgehb3NuXKdNP7dArDOX8z4EX3Hvk5bBv4P/syEkYXzUv+mtzVBwd74x1puK582I4N9
Qlm3IrxRO6VQvkggghqzh6dVG5dPm3zqusszS9d7HoXPjaifXRJlLRGM5DwMEHeCWJ0LzoCZZciF
JJuB9Q/Rci5ZKp7npZUSJ0vLV70AVzli9PKaGX5zWB0smjBqNJ+bQAskkn3Z+WMcRW3m7g36acj/
dP/gYoxjAL3kYUjd3mj8Vaqn8VoWEyGkpyo3vXuSThs8FbmZClBnWr53V14aJYDxqbI2EI8rz8rn
5WiFYcflQ++rYj/4h67h1D/JW+e265NL0o9eS65pN6JySCB16mnZzD17DDf3GIbSe63BKwg0h/y4
nMoJohnyNILj9wUICthcGXyshGwkTC1/+Vtt00OxJrMQwACDQge7OhpLurGPxaO38bs0jW3RgwCd
VpEZFvBYN69/j5n8qQGkcdyWIr1DoGsbVclzPVfLC8kRGtRt1o+DD6MI6qKZmtlTE7Z2WJb49I+3
im/sN6gdT9ECLzm1sAv1aPjdxHU9b4g/gPT7SdiiF84jQ0kGas8K9xHI1Jwo/lIv3aDS+d5PqDdU
73DN7w7HmyFVE2BGY9s6EjH/WxGq3EWTMXJFpM1fPnyGDCV5y12e0Pc+xjMQINR0PVqFqK3YrM/o
4nJA2t7Ai51R5CgBts4APOwd8gXUejh73ivQfTUJB2DgAEqnOmlxfauD4ZOSeyObWmbIq0J2EMwd
PYWxJvrnJH37pAsGloNFLi409XPQzP/o3ZJhad+segNDTz2wxvA/IkWWnqi2Wb79Gpm0A1hdErYt
CczwLFr4yuBfzkMSyUFqg4DrHNguWDcxNhgbdeSENsJCHbpzu75ZlAQGqn2maSm1TlRUtI4S7uz1
cUxr8QnUu1IEGCu0dyXfSglR5IL0XM+JqRP+issPhlBTEgzRDLQX6XYuyrAc7Ik0JfdPwu/bfLqQ
2Nv1c28ItifEI1VIq0PSMn+GH4Pk++tP5rPSFqRY4ZuMtRtPyzsWjb7shFyiEzY5cnZ9c4R5h5nZ
TwZ4I4DKEMztbUHEXTL7puv8JHb7l2CbFQLfqNrjTERvBK/p0GD093hZJrvffNsqPja1Tt28N0Pa
flDoHdi24x0nKZsICr4iyhfenbOYxzcHcbYx0/jxi9KD4aFvijqnpd/S4LO3e9TcaadiRxZ1QsBj
0EXOHNCgOGoyGFyxFpWn0e7LCuvyB8WqgTKj7uIFxmB89lsqTwo88i4QgCdT4zS9W4g5YA4853oG
ZqK6W37oyZfPbPL1kclUAbiY3bHvpXTDrev9darp0dOr06yqH9uP98lPeEnOqCkDCxu7KPC7rXTy
FIkR8Tt8k45Cz5EevgaTIKzvCA+NW/kjGj0X3LyDXhINEiZefv4S8CxfcBJw+HLGnGcoDi1kalRw
1c5MIQU5nUbdRAvFZjNuZ0YEMvgtCRr03nopSM7hF9EGgfJgdETiGPkSR52qqxylmKoY2TXsvIZD
A57I+3L9KSPXTmv5+0VZICiRz1Lyf3THDY3jMqn3oUFUYi3gj5cgcuAIhWVsGVOLvYZ6v+fYTyFI
PXZh/PkoUQn6PJRGPCj7Q81ASzGZfvDwsXtiiM0OqVq27+zIAe8sdbQtg0kXjw/A8qdsTcHirmcy
kKKzmKS0Kr2ib4fl4zwEucK0qyFNrQuX3PHzdpvyPeSKJHfxYR70GhjE6HnkKhxYqtAsCObJ4FJ+
IVVEuAoQUsHlIDVkxkGfx2NmnqxtTYGLqccebPxYgd2mLNsQmvKmQ4J/7vEc+GIg8TI49+iorpB/
AA3Or2Rekt/o0AhbsdATFuUb1bJUmPVuIEN896vA/XX/a88gyDHoyy8vDdR7rpQ+fTie8BC3pVPJ
9EPP01Nqcd27dmv86rY95APixE0gXvq6i8bYkZV5axS7lO/2QagZn4qHWugtkA3Wb/DhOkMCv2nM
wbQNnlu+ujzcX5QYw2ml8THim8olVH1cIC1930g9DM+DmG+Wf5xj53WtzAzR/IGjh8hTjxCSTu/4
4z7LGG/emc+06CsSBH7fhcVXM0XoSSmKeeiHZon8MDep4HKy4jWxv6ZWCfGOjcyeT9USVRNtFo5D
XChtyOQjAlx9tBvfCTmmvD3gs9+QvWnj+M341pBdok213EckJU9Hykp8arvAWF36nL+7KMjYIKb7
xwwB1p9heO68QZDNn03UbkPqtxp1KsiwNevMGjWmFLR9O5iCWJ0fq7nilcV1i9+Q3ixzdXpsxGOb
jUAcGn8fHkopnGXSWUIz2UkpXhErGCIIiFVrsehRSE6c66A5AaOp6oYUWkHuEGLFv2mxN4OSxndW
gghiQwkxiqH5i5pkOXR0Pb87LYu3BrFEV6Y1VGAAfBvFuXxpg465UqFFAUcjVOOSNZyxvBqKbbNH
c55xsSDnehQJddyPeEbi2/wnm5QrFycIbVPKhU301Jui5N46CTvOmJvAHJ0zWnr1j/32IlgeoppH
VseqzcRvgMFNxSk+3MNTFs2ZaaAzaNU1XIo0Hfnvscz9ZS2gnlkAKGYmKdR50vWt6Nk+UhKeT9nB
dr+CMKeq6Dch/dE9akrN2EJzM0DMPv3Piy5JG9YTTXkagzJtwbxRDnzJE5Erdb1GpDC1+SXUn7Ah
XoLb+6XzGw9UtqOpkJ3tTv1OKqbCZwzZfRhfK7HngRYDcSSqSZu5azIlMh+vnBZX6tWSK32XgHdi
EuX1QIKX0JjenOcPx/Ke7kvJ2djutLKq0q6iImC1FnqtrtSxssxrAhu5Xl7BnqS3gf9955M+6P7N
RDpIO+sbSXpSyap01+BXrVeaGZh8HOIcJG6r0uSsWhaBnuRQNbi5XteYHdnhcn4u4Ya7g3pDJLYC
ojzsqAe3326feGjBykJXoBamKaQXwt1QHnLnketkv8Pw2SCo7q/bClCfmZtBvCUiA+c9A98UWddi
AUyPGZWjK9R1Wm/5/a2DiLtgzqeDujHNoHqVixIggB3xg/bn00iLbrDuzR8KM2q4aL4gi+A0Rr0F
OrK1SXTFrZPw52T6qV9Ni5GRPT1RFJt+cvtUtbGr1WqrlyMkMAQbO/nWeKqW+O7MO+X+fksMlYMa
oKlAwUuG6mL4OrkdxeGfYPSKnWnO/6t3kdH3LFWxXUwKMNnV9s7jS8m2pRzlUlOTDd3ymx4X6mK3
tF0j/NGk7afYgQZ25tupqA4PC8+sIhOU21/nrCuafUqm2IROyhJ2EnBlYvKsW1xnKqd4yvcr3n0C
tjXejnvQrbSzkyz+DzJJvjVELG0Jl8DU0rTBy/MUox9LSW+V8hB50dQsK17v8MtYER4oo6aEZM13
4zSv1gLH4RcnoeyFL20cuhV7w+wWMrsegYiI5n8gFIZyBUdpxsf8cZVwxIzAA4cD+EYg3wnudOs5
0BbkhHGmqGme2DQdSdiZ6CrS9DS8ArV/xFsezbDvAEYdOPlNpBNRLk7X6B9H/dJ16A8yMkXDjqK4
YJB1JI2qCEa2Smb+p1Xx6perM3guYoMBH4RruGsNOSgy/AETf1aQtIr4ojZfFs0bQ9BgEfjkjrfA
Oq/8j/t5SQgxIhsRDnYJqr1HafLdj3o21ecaFSVBLl8oLQ8zsA7/T2lT4gqpS6sQHyxME2TGaeFt
LxlDrpOVOfFFKlzzD4ppGcq/89BA9L+wmcD4OwfBlAmXr+HzAc/+xkHox9vdM8j8y0IyETQyvGjJ
pGItov49bWAmS/vsGF8MNfx9ednzIdH0IqisXVaqsdiFeumnu83vCTkfOSjrzWD3MacmduysP6a8
U6r7N8I9fQ8EkBG2oDPGQQElIPpVe1eCVT0yh0JMVyEiAryHsh8VbD4Lj4BPDhi8dMgJfQkqeRHS
4nrU9R5UuoruBaSR9X/bTO+TmHxef04aam9hC0XgfVJ2T1DfO01bKoOUE/qw6tMMNtv+EDEpD/c6
e0bCOjaRLXd46WYfnjrrx1d+y20k1UpFaHpJTxLTB1ewLcWc3ezdovTpK6RuwqouiNqFw2fXkHYs
SfBXvnNA3hGkUE2OU6hQp9b0hgudVRDCSfNpFgk6VSmI8jnvIS1YtYwP7Krcano7hJc4ZM93CaRa
jFHk6utz8lHAkbkEqAzQwas40pidsNm8ZpYXE6PX8ve4psXoWK5X9oJXmgK66NvhmLtTgeh3NK2w
JkFYIlYnYeI5cNVCdjZmVVMUWQYVix8k4XdpORQWx3HmKzNFX3Hs8sYrgjVVkXYa2NQGWyQZhjFG
72CbFSpMxrh8O4wc4ZLEFDRcNi4RcXaSa18Fz29bVVbt6ysfEvl1ixyclYFN8jw3AQo4t8Cb9lPf
7hzjcOFPClIoc9WPnzJJMZaYeqFA/OiYf6S4gDXXinBv9mnRwdz2gf3cXMyHJIWXT5aBy9hFOu34
JurtmV6BLh/1Upwlwgtl1lLrK3lGyYAOcMwdmxB18ZBAZ2wx7RQeCLjvbqND1dOc3Ummfg9at2B1
So/EwE3EMYDly2t15GcViYaufq4oY5o+EF4axhBjw72PtVtVjy1BOK5CKeyXcWsWtccMsJ8aF5W6
Lt6Z+BqgdapIFihRtJOy9FXWsQjv4fZRwC/j9UTywYzU3Pvs1G4Z9OtDNgNpU4TMbq6wyeli7uym
ASvafID9Egcbuxq/NQwFVZjiWtJr+uGcKe/8P62dq2BvkDO9MEurXzm0bvjaFLOSM74utopyVmsA
zUsPKciraAmWVG4j17JOkmSTKNNHnaLOxSjawkH/LXzBWwN1fIFcoGEXa2BHHd3ER7vRsePcQq3x
1Z0Evadd1YhH9j48xNoZ6+/idBj15FxD4KR+L0F1i3MtVhc6BAWF3ztFSkUURMv6X9YfPE8rUa8l
F2gyRH3OQIzX/p8+97yiaBiqLnkYC01qMK7yMOw+I2eDdTL5NGElqVL8EGnsa0SC9j9YYuUGh6et
4gyusNHlXm7zxNs+7CtGSTt8y43Uy3kFK1z41j0xqHLyxe0BSFOSb0Mq6i0MTRodF+oFnMkSd4gi
Xlob2l6qQFHOdfVH91jCUrh+KTWPvzUnCpyok269kGR3EwjIxBgOtiLYWcOVWOUjcyAp3vAd6qGX
Fxaqe4xboWBdZRASGHxh2nc3SByXiEUQ5lf6FQW4MN+f3QXIxyY5GiqJmZQp5Hvbv5zHTPgROew2
CG90SiXqJyWV+Bq8wNJcpQpNzd3I3dULwjI+2wRvmvrO//tXka9VzcbhG34XYuXdinlq4IMDqNxy
bN16+9i+XPtioo/ON9uETuCYjLXufRyNvjXhd4/QCF/CwgdzQW6SYzWHCk+y/x6O3bqFdPTddcxK
Y2EvkytVu38X/Vm6BI92mu83ItI2hDtcCZb988IJqeKpkIkTyqE0+biMouSt1jvUb4QnAxvKNdVe
Jg+HiiBTmYBIHc8fmXYZBCzCocnlaN62XdnJG1+20Q+HHuL6LaIy+7cFZCIVk344Hxl4g2AVLcv7
JDR0gItyk0lrFLTrp1vYzWW+nO6e0G4LWEn+6XqCWh90/BUOAJI/A4AY0W3jKGI4woeLE1VlLEfd
lwpV7+/LrkXEHtT7fc66idzcXZybg2T/wLM4UqvFIlOk0D7Rzb7tlwVt4cphhFuT/KOTUxrYph4O
eFgsPZS9y2GVcyUl08swOXXzEi66lfQd0ZcIGdBpiP2MA8m/apSqcEle+AR0zypcSYBn5NSOMdvQ
bJDSzxmFPAQHLhe5ilciC/Vd7/F498hZgPxk6YA9z04gg8H7rbdeJsr0Co555b9tFV9wHDQYYGDR
OJ6bJnKQh8hD2Fu6OuuRgv2uFm6cgyBRcwaugp4sc6LlLd5tDt5EV/WaM5iHZJKGkyDsprM5fPaD
MW25pgUspvqGSuO5aRriPLkDgID8HJCqZzlzCRbKR2+5JvJliHo4BPv26bH+RDpvN9TJ7X8kEHzq
I1xfqXxrYotac8l1JCDqmi1RzX0UE92Ht2jhceEtVn+wvGyLaHhz2A7Nxt6oOWhpPFKtretlIL/T
pvBgFnThck32n4Pn37yBdnc9oC01nPOJdFXHJmZADPyXeycBN3tDagKvREPLmPyJr+kcqJjIqy1T
+Pyq514+LaNs3qBxuDtcajVvE61qAGAysDfD4cGbFFaF5/WYcB2RCqMenWQtHAQdBo0EBEGjygfS
kPIKio6YZzr8vnuvjBqq4yUw/5fkgMT7Xmo7x44klZnwaWEt22Y8tTk56yY0QDbBnp6CHrBDwiPH
0A6EE3Ku4cNlDzgWYP6PBqrT9MLQiyIl44N+kIv75NeAxvG61gRVx+cmsrLVndmNpGxjU4Sdmvx5
QMGXmKbhdJaC0ZCdo7q19n9iEWCACqL7+JrDjS87bcAE4biUo0/5fDflPkyQGs9DBl+KEL57tZRx
VK0naXvenW9HA4eoKz2qTwpnqYS73CsQw8+AYodCEE8UXa7jGJjhnHZHDGPFojBdI05uXWGW1J/3
k3kdkDtz6uqmiKFHsOPw74jgfs30wEpldMrsOfcRxUKH6eKkNgV2XNnj/ba8suc13tIJM/378/ak
LYaCz6Q2F6/UtHpT3nR+MAxzA0NxjZR3B7OwOQYpCwP5gdJUfuDXaUHBGlxx4AgEDGMHCjVrGcEY
BM/lLVnY1Ck63QpqJAE5+54ieHRRR9shbj8YGDfTumOfoCY68Zc124aoTtLYrTpoz6uYxvwHPm5i
x17gFJJNCCGfSo6sXMM9VWagHfAHqGI2piVm5PPOR3KlbeJv9UcHEDfW+seGjn/4UnIvzLyphs/Y
uYE8qg7V87VFODgbXd6t4SXx7qmPvLBgIAQsBKhUWdNhsdD8AwVMiqu38cF6/LcJhBbKZoXK8ech
CMgFmdy73Ne1HKNnNn6MQkG+SFv8QS1MwYZ5k8YeMnc9HZi5rswCd4cxTHylGfGDtqXXKcWeqUEN
KMxNx4z8asTI042P04l5yC//Lbg+Pl7dxaQLzuI91CeaGhLbbhhAGivtuHI8P6loBzf7SWkBK+fE
/SQ1ycy/J6eBUELn9cn+vkMmnpgchVtC4RB/nEMPQh8h/K0QFlIIpamp7Kv69vw6iV9UxPCoqIyz
koCsNMq7BjNdN4H/07SUmBEmWiWz4AWu3mISGDn9I3Ne4K+fQpOlssfqyhc+YLDBAbQ/oGP0rTaL
yxRKlYGEDK0F13GYfBzlWbzBdJ1sfle8h+5NWC/sEtr2F5WTLe3DYhmz2eD0iSonbRCvefpxpLTv
3G+Q62UarN0yXOhc5d9/kGYRjFb0AP27r20sePwHr2GYnONv8gGHlET/iLHcrGU23lAGEHPdFg5h
tjQvo1cu6dFCx6S2dFu8cOR3CEUWpOdxw/LfpZ6MK5+RnurKDq/asCsV2rh0lEHwl6FH0EOtjjhs
gnNckNjDM4d1m9vX3MsRGoIP4yOuadyJXag+qDSWMCGd12CTBkpIQeb+LO3r4UL31xFw2o02gvQa
6eIr1ShUgt/tzf55/7Oh6Cgd4ysCvz0eGDXM5kyJ1OX3375Vvv7EFmR5cFIjotkWw4kjeyE0hLNR
axD1m0ZRshdTYo4HLB6FXetEp3/gPAvQ9dLuYwNMZoGfeOLReBZjyeXJ1IRowpSJdCFKfjmJ1HCv
HirSKQ3ratBGXc8GoTuZ/3DGkJ02f/q/sbWVWYlUlFfZEZ5npk1gZXe/hblBywifdLoleHNCUOy4
Qka/8WOdflPw7NfuN09Ds8Bw8sO5Gmy9xLDS9/fGgT3rphWDDAgO32tapeSDRmcR3ahIJkfnGpJQ
ZcUErsXT1z7oUVQnsl82Ifnt9AvxKRjcGaqO31r5Ozb+XP1nnFFlmVZcd0vtosOk+flObN4SP7k7
vSI56kRvcUwfHV9ehcW1yUBGADlr/i72SEy+4GG4LNwXOD1Vjm3av65OlwAuQYDpAFtPUmTSzRbG
f7f6fBWYgFGqQEJhn3gd4xJ3jA7UrwDEGzgxHGbzK/GJoFoXblgIQg/uoMRXTABRGLv4CS8Qzu5s
rM2AuX+e1RWBxZZRNXk34ZEpcbOsUIrS9kbqV3uHDLvweCFcBy7IkTmqn7uwx0qgKMOZ3TBdVdxe
ALkz950ok4VUCHqB3L+7/ufKY3AKH/8LZqqARi2hLuPq7mVk9qAwbkr1ztjHXRiIRSQmBDKGgK3d
VZxslfs5gvpCVOd5E3AqfBaRNpsbBfWgtPC26KwoItop5vHSq43Hl5mp33znoqoER7DoxZKwDpQb
oTpBSSsCPXaMWxu7fBBsdnTjQ7SVDxLaR2s+6IS03q5uk8RNrq+Xynv5l1iw95yQoJnmTQfN7xRz
CKOHHCjPrcA4CFd3pWiR41N2TOOLsgMWgnFiOVAu2yxfuv9LClUsIePRZ4sXS1Yh64PdQ7K+nnn4
AjcWhJIUfMsb6B0LMlbhTTktTCojdCJOlYQJALWoZwpY7J5cn1tmZ84VgR1J8jAC1ByEK4Tfm71N
oKX+p4wnw3Jt3MokwgSUz5zbeZ0K2Pvw1TeSvk2fOIO9c/acVgQlnQAqLdvDcwvyKApoWf6WOR0U
Wnsm3Jv/pWI5sjzxK7iZXtZWLFob1mhVyL3+eGqhObbk4WwDHiXiwuzV/idVRzAJQ+ttljv6A1Rh
RjmDP0XXuW2/nbsZxYRdAUFsmaDN9tPHBS20FinLitfXWZ9hIJlTbuPpwY+zOnPh3IhxmpAP7rma
SUFX/ZcNT+khQGPMiA2ALDIrnXUcRL/C+ehpPehODzJwg34AeVBJSHHhm55sJK0ZnSB8L+8IZjmv
rZEji4mPdMg4/4v0F67FFev+p00xJGcTIVp4L6JTPIj18R5xSJNWLy/qbjdql1mWycNyrlLL8Cah
eAKRRkdMNteXY/FaTbE1UgvaPCMSmvk530xamw4VUJj7b1/rtm88zR9Ir/sQXN8+ID1RNhAbPrVu
CRGxYdq46tDdUF7FPESbi6abU7XAX0tfh+sQJ8pqxB5/Zw56QhWjvyjwdqzgYg5jvXPpscOQu0wY
ExA9MSAXbECvWRz51kxGtu4UBZfXpVc/AjglYwPiH5v1yl9QWB9qdnWrgmKAbmY6DctwnwEhmAIM
KI+0OKa50MSd0mwV9jBGIziPiMQEKF0Xu1jfZllmovxmy1Eh5Vss87fMe4J49Me7cnh1G0xCUCEu
7JzZtbc/biwGI1/pJ3nL0QKLxrUOYKmgq5WK8Ntx0c8zvrRjvXSNVGH/JDrGcN5FyJ77OjRht4VF
s4Iigi0+Ks1RWdu5bSy1pGg5ywCKyZjI24/bQ6zwYn1oFJiAsynWq54dOAhgEOGZu/7a8at6R4p1
Q7VKcfCmmIoZw5HhI+IuMZozameAJc28JlT92iMSldjwzYBMsQzprSiqa4YwRnvzEwA+epB6rywZ
9RV6AuSAOV3riARpOAvdTnpLBo8lfDhYE+xKWqje68JbAx8a5OR0fYrD2kVjkhRg4lMr5OpD1uaC
LbWAqDxUN1ee3hsjTInDkymkRp1YI6FIkN6HPGUI64dy9NN8qqnxWW+emuuZx27ChkfAqfD7lDni
kZQF3NSH5bfE8j+5n5L7SblDbLblyIY15a4Kmn8hI+7Z0HAvPCctcgjrMxkresUXZrf3Z4JZgu1F
VNDwMMCTCAAPKiGGRi70qAreyJgGeKJTwsehmDSPP/4UUsbD8UjJzXtJ3SeyafSrjHIQrm4WmKKn
pFHLC8wbS4wM8WD/7/cT3246lUzE9hsgXckOSSBgMNfcf28A4oFwWs3C2J/Hhtw62sj+LjzZ+VSh
3PPPao9dX5mCk9az4CG+rP1EadA1nVhnsJ7KMtbAXas9w62JSGb4Gc+M6/gR6ywjG39edeCQoMU0
GWjCslHE6HkO1fq7ZW+1ij7H4PglHIA1LEuzWsn25mNKWPpwVpsw6kQtGKi1WAPT4ZGEUd4ugavr
yIpdc9zHgIUaOORCpPDYznUvYkv1lsEYAM5Aq5jnTbfokhNYkTw7d2HifS1VKUWN2s8ciNZNyu20
sxuFqkwDurmCDpWnU7S7CgYAqGs8EleMDmgNGwAd3wOgmpZodXUn4KzC2iFD2yiU95WEvKjhAXlA
d+5PxeKO5neHEBQzRRRoWgLXV/O2fxJ16JH2PCnozXvOhwBZidpjbXNLW94PJzGujsKrAWSjqpjB
EzTd6C6PlR6DWHZOsClZcxYnig5WkCiQRK/79kiX1vjUhV+h99Spfm4rB9sL6EwnVBhkcxW1YN18
iR4vE/e8U1To0TiaJGym3fxJhlqoZ0sqLKdUhspGu/uBWFGeRgwzGDUIiWChZDkiTxl/O6+fT0AQ
Iz9WdMxixE4KXga/rMZYunbbFG5ptqcknC7I57s87rUHELVfIGnqqPtlS83o25qSIAbg6fZ/nCYZ
4NUIud682V9fecTWfw9rS0arEZA9WVefDjJGQKwe5uo8EWdgAnLavrrgTJ68Zt7vN8+5uBNKHlW9
cSVdEBJabAIOumEf2f5vqPEIVSFcuZU7YgjQx7DRFCw1bJzlt/4OW600ydj9M2n9qHan/cVoYrzu
4UE7w9hoB2oS6GuGieNkX0C13Dudc10Veeo6kEqYKxHVTwyuk5r6RAhFR9wxLEIaPPS2Uuwbqti0
09I32QctcM+2WCcYszH2JzLpFXZJaYjNeuA50QW79H3uR9k1+JfNRtEFxChezEDwIYr8u2HYM43D
5tb5t+6qfkCbIO+jDWCTa3kbdvb6qRq1APEtaml2IpVGlK+lLlzng5IOpBerhYnN+c+lKylmhJSw
p7vPpkGu4bXy3AAKkfXb8dYi4iS735bhnp7ouw+kLWhtcX3tSA2vd56D0BrAxqPLb6F48xRf6sCs
FkBgOI/oJOHXDKN2/LIxcDk8D8iJUL/tFPWkLa1Stb94NF8PH9oUDys1UtCC6Wc0C/cGKdX8cuFi
6GLmymkR8HnGMsG5cuSxkMxQ4G9sRRtJ5Um6Dy3U5O/ecDqFEVY3ZuyWb0v+KAcz8ppUEL5KC3Sm
TM3AsZ0UcFUD8bMG0+ICojrd412dmZ7TN+m0qGyb8b2eYBt5CWEB/mYxUv5wvhwa+5cgV6GK7QRt
RIxXH8lAWQY9wbT/AMt6izpjtXfUpO09SWUf5jw1/4tI4rD0qkv1fP1UApN6at7HFjHfDNfCXpp/
9Mc3tEpUV/D3GUTm1Ts+G2FH153DCwgA0YqCZTAEgDcN49E30pafL3YwCXqTTPAObnNo2u44pCYo
kuxWl9zWsCrMgD4bZ/b979kOJWhLHrxiDMxYfWFU/FK5kAFZ/+AoEcWG/WxXNJcAIvtiUBwQhneC
UJ1mQa+S4KPEgDNsJ84unEfIOoGXjI0EBnNXF0I0ZJIlyKKDAHoqX20zvsSo8o11sSAod9sHOqrk
8KClQYH4Jt0KbXNO4nwJwqr4Kzg5WFHx56E6m5VvgpqMDegK+xMKBridIm5eEG1QTuweqMR/UspS
Oe+B0coU5FGRWQDmvdghUmyASF2EH+OXXcJx2/Z0oDljHdAbGkzShIVVDEkJFWzHa0cB4FsA1qKg
cRK1hNv9tCScbTrnQGu1TaX4jpcByev+1VgzEkWKX15VhOGmbHO6T/A9tdAbLd1qcxvCr/yngJQR
xSgTaK19G2tGmhw6Fl/mC8uvbQXkcT5HiInlUdD7OyGLlz2NFRgIXI6Kr2iLzgq/LpVHJNLAXhy8
kb/d4H6T5cOQLqBwPikNugFxv7bjvnhlj5tI3/KS9Mc18VaFiXbLKr3enfawPwsVAvNgaoOknmZA
E1BT1Xw8d9sOxkR/5CUji1E1FzsdIwDRBzTEb34yPkhoawFmWGjPV356WIcJD/FDnXpQ3Bovwfd1
TtESJWL+sr0ykNnRWMuN3EFTUN2HyX1VWfv1FaxO6EL2Uk43Ykc0FMabbGHSLnTpNUfNmcH2pq5o
Qm7RFaBK95zOwNQWz//A/w2cMdA30MF0HL7uGjREw/FruaE3wvFezu+7GDKqMT1TIysH+HmFszE+
16nsu4xWsw9634iEt+Hf+Ty+7cB02q+b4r4WAu7i/p9iku0mkOO9uUkxzctXa+0fNMnwVN7+6NIk
m6G4jsd6B2W6WzbmZl6GOS3GjFpWErkvjVzyfVgKT83LeJZZa5XW5mlw2UZoB6kj5IStViOi9DfK
o9gQPyca9WanIX5MtP6tSp24J5QvhVMgPw5Zok2kl1xIMaqKP3/IikZVRCQO/U0NLB3oa/VlMrvS
WQCZfLL2qsXxk+3pYoWAP055XAAzKebh4Go02U+0oU+sfP90IMhG42Tr02bM4GHut9LgmgHCudVU
67MvrcklCRqg/I9Ad2WxkOLoY9E+Hf8aJbeDKgwu5ZdO8J+5BwaGXJQ9CKETHDIROMct+a2KqwEd
r0Rb9aIa8pWHZ0l4ugrcr1zn1FyxlV72luaQKAxFhN56K6zneS5Hj/YK++MkWlC/k+xZtWcHQ53X
6oRAMllWZUO+dLm3TZCc1QZv9ncUQggH74YG14KJOOjqa8GytRIf+4ytqwnhWAg6DuIwVkeBN+fG
iARKv/OVnIumI9/Px7YKj+eLzj4n/KctPhpezoMWbwXkzyneXiDAJOTUA9ZlEq62mJg1qnL5ZB9E
Do6/p+Q6yJS02w6as4VG8j5vf+LTBgGuybIF9SJ1ne9utC49G0v3Sxd5ob4MX/c8U32f5XjwehY9
WD8yH6UakquGQwWn7OMvhmQuWJIolwBj4Crfn6kKUcHAhqjMCituOP59YvYowUXAMvOG/35gZBrz
YwcZ5MMQNguSridg89E2MYz2pyqmDSJmLHKx0GGybX+pxSCIJHygCe57m3ad1SfabQOAHlXaTymg
lF+c0PkaelW9bt3FEJBqI+g4k+9/d4CDOhXZvyQqoT35KwMYlFKAS7W924Xzuy3486kGVeii6etg
DSGjIL9BuFuEZt/Uf0Uqv4Sg8SOk2WF7fisMRHEbRxBNyEzSUZAGA6HweUjQntdeGK5k91eG8Lv8
wAOBc+Lx1b3lK9SjiZOAfoNxiu7CyMHqvKcQWcul8OEF7ZVBRYXmjZMMH063SRaV6F3SXrH6HF8B
xhna7zfL26DVvnclGRm2fkvcSP0RQISEvK/iLZmkA1IONiABmR05rOA5bxk8yj0R+oBpZ/f5eZdH
r40hym/mcRkHe4lWnqEnFXauTN61NMF8znQa4TRSSN4yir0v4SgI1QLJhpYZBKKeDxaMVpazHfdd
UzGaJRFN2CDzTUy4PnF+NAV4iUMyrYESMkV2ue7rPzyVZ6aY8doX+8KA6MY0aQfxZpn3ITo9t4PB
4N3W/7ygCXArXtTZm8TSZhYmvgW5fsLi1zqgbMm/4z6zsl7vNhgPHy4HkOf4HX4db+vo5fp/g39B
9FXB5D9qbOg5WERrpjD+sdzhUDLEkemlGWDV8HHZ0jm1EMwDpy/tltNmyB+y+nNoqd1O/3LFbvmy
VS/wzI+A2s1f2VI0UiCRT41Uy6vh31pBmdYCaEvSLOtQ1ngPJEfCTuk3C8Vh6zX48RhxrQciDAqq
73Vhow9AavKPAJ18xWJhBOtslR4bCjHSWHgJesOfPYFL+tP7uki4aF3FGiuXjInBLeymcpziUdNy
XjfGskQn/fDw1H4isF4KoXk6d0Zabfi97WgwPP9F6bvWBBbFYjKac6ozvpydNY/2hd5VjzaJ4lzi
moY+khJSYNIKPoTgS2GgOsM3PU3hQfIeAhXGhZTU+Ta9sSTIm+fggLpVxk/gds+9tudsGt0OAVey
gbO8XpSryO+0lNOeqAuzqi73/v4i0+iqQasGJVHovpD/NuBSfxOapDhqQ4MsPjzGe2Jo3KQFa8a5
eidq9GeOo11rSV6ydzzGv+IDAOcAo1hL5KHcIdjWMCUgXgFy2IMkAmffsmPndikot7TdwyGMxlxX
c8Hi4sbJ9wZhmkjwuQJx2IpOMtuIgcNcUuedPfRHjIj5qlLtv9Hc8VkDnxI/6sQy7N52K7gDIdwJ
HVJ6yg9kR6UX5wlR7kO93ToTlTj56Qnl8bvbnD53dCASdsyx1umdRLjHgciZpeaeO5fUEetMAEQt
THw3oNVOGe8NqtNiD52F5XW9Og+y0kqn1XttrHePE5WwbHTiU5AnAbm5VzmeMOZR9CxVhHAhJE5Q
gM7mfeKzw9EXTcCunQtco/w6J2aNOcGQ24y5QqYkAWTa4J8X5uN1pJy71/LrwhgMKAeLQpU8CH4l
h3ZkfRKKyG2ZQSYh8+tHpwwQXELdF+T7cQngqr4NjSBSkv3In9tKGjbUqocwK6twoLPPVZ0SRp4X
SKL/LJyrqjTeh4O3Boq2p++Bvv+rpHO6XGuHz/tGWpc5HJBE079KOdz7WIV0/VFMfsunX189NzWn
qRzUtXfOZvIMKmDiMP/IIvdBHAsBVu5OMTCzNaHnNMrRfJG2tA5G8+UB07pNFaHs7pskFe3RGPDS
H1hqz6R+GIIDd4ugSqELYPLNqY3FLssn/g6OKrl3S6HXOHNzn8cm98MSyLvR8i91o6xXl6d1IaGx
gu1n5Agc5/AfVelye30p7Qg0UFp9J+W3aWtIZgzGH0qgU/kvHK6YUgi/LxCu7z4U4b7HRVytGfZW
pzmD7UH4N2CLdXDkDD2dRJmxHw4R1ZEwBBqcCZ6zHniCx8a7bnYgWpeC4f5lfuvN4ssaaVv0IjRu
FhDyW14/q95SQStSUC0btm9zsC7IRSE5GjpCDSJ0nbeORKMi0vLQr1ML7oB1/Q2+Ow+d9SVK3lhC
lPjh6/SyFOqjYe61y0TQ+0xzmOcxUJ3vRZx6mIre2GqNNGl+i5hWcvTJnF7y4K6nrJL4VvUVqz2c
vNePVNT0Xa/FW+lGiKdfuK8VFsbB2n/5Vd4+7kzd69rFOlFhs+A5XoDWlzOZDwkYqzDg/3+PmFzH
ST4e/RlY9cNGlMg390KuOZr5vf/hqTn6xbDVgsf7wFSsQT+AQNs7xkIgmdHAtcBnGfi47bHPjMth
r2GOHTqooNrzXUPrmmJKii7pGQPKNJEU5eSYTmXeNxnkvKNJN18f+Hr98zgS4goQEhTL2EYQFXw/
MfQeqAttvblrhgivSQbQOnMd2NJtaMSDbuCwc2xeMM2jkznC054kwIeQT+JSA7AVbGwd8rxgPCYv
nGXf4P5DT3J5MSE7SsVNU8Hlhsa89wthXTHnax6Wnp9kIKCjfBC+MDKXQnCnxE9Iu2DvTsK/WX3o
Ulsy/5asd3YwTcv7ddy4A7fIImcPllDHM3MCJW2GgjQ8/SZRAysAWdWMK5qdyeVgSVNzehBhsLCJ
kh7xEC4DQ18NzsdBwrmuPwOWsdMd42wAObIN55bOIU2/Z7L4lA/rCCrPmCETCKZqUGJCBPRgA9Rm
c9ZV+tS40ZwN3bI55p1E4o0h2QAnTZJT3S/V/z8gGINt92R7vGzWkMFdzx/eu59i/+gkhomXwdnv
GXxPDUZehtc4zR9OLgAnFMnSNRZpwH+km1dBqNQ3+pvsGdgsVQ09bPBvvFVxz55Ilo2XcO1Kbv6B
BquW8bjApHAbFh3khOUZN4yQQ9D46WfSFu7d9wEVlUKZ83AwsQ2qfd3k3UtMV5UF2gcV/F7nX2Kj
nlOJnoyRQUTWJBx7ejUi+MXnLYElgNG6HazdvXSUq/cyyPMN9eD9q4XwEu1nkDH5+POLoh0zZf7h
CXMYsarK8/LlEVKn7vayPl3HVTHFBmawG33/PjgFM1U22WTHQIxp4uVMAEan1sC5q059iSD06sdP
NKRHYA7DLee/YhRm6BohCRX1OcV2XAoPXRAbKsUGlm66LUDcg2Te3qBqJaKK/FQipmYyywa0MpK3
zx7TDe7pKo/32NzWygUv3eza8Su4+NgOouE715C92H3Ew+3ccameMG+AsCqoBfxDd1ZIWPKq93+M
QvdjgjR7M+IxOyrCUBKNtC0uRXsKe7JXji7FwjzKkE6miZLvGKPHwVaiB276bmiRy5kFn0h0Xemv
xupJQsAMyYRLGtvWQGzef0c547plCZ+QKl13ev/sKlgldiVP3bd1M0VqEWJtq7ybt8IKcqGdgfrW
G/7XMFbGI0NoCXEwAWWUsg01cRcdfsjKGgUkkpCzZs9C+WjkQX88gG+5DksS06UhSOqSsXCWO2C4
7LDqxVEsdIYHk4ZnhGyY7M417ReAlJZ9EsSPKMDnWrG6VQx5ZtV/ZJrR/hjv082Vm6m5oov2jGY4
hnvfRZjRn7PK5J+Rg9DiG9thYX1TK+N8w6c6KTdOA8jAraU4yoYtdaBe6zvpp+5mu5iFoJvOWbNl
AIeutGL7w12PQQHRtqoELCe71svrMUEvZLVqA08Dxl2VTPI2lyjAXTpHoLAKQxjw9N4ovDMFlXEA
TyDd0clUhKJl7MyZwsynQxq7UeF1cdav/utA2p5AYtHs+/6Sve6DIfaDnhxrJEAUUzFtnK0T+BCA
JfdThgHVG9e00b6bdKX3E/evsdTjwNL4F6GmTGsRVLHQCJQj7cUEpwQ6WCzkFmduZgG6YXteozdm
2s9jz8iqwAkwxLhAeHX2p5ma5pOE+iSnOv4a4MUzOaA6khb56bZI5oHadQTTDtIIgZGNIsvzrw4o
7LepHR2YHRkTTQTlhk+1oD95q1kELublGCvIhUbIRf9G9a4uQxxWg80+b7AT/U7QQxCOrcOMKbWL
S3jVZufLrYWPaNDQkd/5DuBEf5fqEiWCqHjBTbe3Nr8BuYxbKazlGvssX0a7yYHy7uolRqUjpQM7
Ia8P35LGU0nxlvcVTC8SvazNYQCs3sxuW3Jg5eHVwpGy8jvEubWoQGWepqi8tvGhxBD/uoop9T5J
TXlhz/ShW5Yx+acM607ZCMBOCVDrXvPFM6jaGohG/++TfOxf6mowCQDQdCRwPj7xUKkNA/q3DVAi
63UpXU3Wu8+UIYXyBis85GjEx3YSKFdElOWA3BzmfdVUbzwrxUNmCp+8PFXRg/rpN1EinOoUd0+c
II2xerXe2YCchK5jP1BGCcdpEC5KJJyomFOctDWZaR6EYUZOdLXbt9bW5RSUjTlGGIIdmAGwXJQl
/Xnt8lVRreWn4FC/aCHRXBpE+B6diCHGqMOzRntD8P7yv9Emj0byBxMIykInpOeyKdqcNOwtIyC5
JvogmV5keks0mgV4K3tBSBn5MOQFBYFvG/yQMXGoSjycuJyUsBLf7ssipgCqUj3JoR6/qW1M/QWi
gtMVpHjXj+ZdRPnfVP9p5Dx8CuR054KM/5UFD3wWbGeUayFyjZb7esuB2G2oW+kZHTVBh5z6rxUE
N3eAX9gBU7Nio/wHK5e7O3i3kwp+xkk14zEn8dug+psuXL+4hY3Mel0w2ycgtsvkDENiKBuT/Wzr
iARMX0Yb9y1RR5SO+OWbilIyJUr5WJjZPtfY1UorsvTbNMBwdDUQm5PRhzYkYfqmfYESkbQ5cqGN
ER+iapflBfC33IEeIKvkveKfZzcdnShgbOqpm4dhIgzj4j79W4Z2/H1vrzWbuPWJ9LpWD1ZnNXKU
8JDVhs50Wjm3ZpPC2V0kCwmiGey4FwKzAjnSFMiSyjbYQchPdTovAag6KQ53iRKMvYpHzGt1yLQm
O1faAlLV+L04cQQ5OnXS6rBXmdNuufXGMagIcqvJ7q0VuNXiCh2DdZwWSDY6FhHeYQLzk+r1tZ5W
/DuhDZxWSPFPiuvuViBkPCMF9v7X54QyqmasYUphtpBg0feskgWQ5y448DhzIR8ysIlGWfhAGRmx
loCIOEUjNKcXQFcvSg/ia7EN1djRVrC79Q6ywx5F51nsSJnQCJTOQwjnwkX6bKXg8y+VUQNSbL+L
4af86Q6jLUL1b1sRXO9nEnIGgaza/jlMB4LfnVhNNSosXOIqRlOMSdihtOXTYxtzw8G5raxb9JsA
dbe1eaBFIvvZLrmYjhII9fr9VR98Kee949BtZNqI8B6b8uuIwUHdYlBmumEDT+Eli0Gk9FEpeYwn
vzH10e41lH+jrLKCxBWWUD0TDj3tRSjJwYYv1SGLP0c5gAeZtDgTM7y4cqa/pUMJx6rCLYwRRVpw
c31EEoUf+89uItGPaOc7s+UcRHu7oqEJz+dDPsmterhQDI+VJXMB93kcrcAarbeP2DgjxfQ8T3xs
RVBeWoWFoScQLgdy7i9I7A936lW+aejx8IwRRK3onO+TcczObg4Qj6b++Bd3qBrHJ+N4GphPmP2S
+Mtl+3tmpj7/N+32bsj+oU7QmADCWrAg5q7oq7EK77BBO//+EG1Oy1smeyAg5SU7oKcAmXFXuP02
qyYJiaVOm0Smtcao4UFL68l2UlVRMR/lQMHXZzailO5WkXjpSV+ILzzG4+HcKRARZLGBbPmx6zEu
FksGCNuTmanbHJUKxg2y8k0o/C8eMXgxX1+rNowUSf3AQ70lqpWQGHoVrChGs71pc9fd0MSBt/Gs
9wVIKMRbPllXuMf+Gl5Te3eZrrpY+gz8PRaDzfAlRtn1Ldxl6yxG8fRl00SdbWMcz5+buCDq2fal
pAu8lOPNrtsOFuZglWiR2lOfij1OyIG8GjzfwIcmYG+ljtV8uKOJCKN/fRWhmJTbgAe14W0d4ZBo
7kB4BUlRH/ZtBP1ccN84WfmYWKwMo3mOxWuAAEpqZiG9QN/la1tEUuDKXqQcq3rdVGcgYpa+w7z7
yUx6xWpnf/Zz588ezcDd0bY1rOGqXr96ijWTObNWalhsV+ahpGRnqGptMiKWtXWFcaFS/SDRuzD4
WZYQM6GiYdkDdJLeQ0+mLmEdFgLw/bZb2/k49tdJwpnOmQumGKWv9fWoWl/URbUPV/7HSvOrM9OJ
mUQrNJgqLX0wPKR9/auct7740udk7znBHDz+Tpv7c7EDFr+TqsiWxkYMCa+JJZNBIcXwJgcLt7IL
juW5tedfkL6pBmOlKGib9gZs37dhb5LFJBvIPDYvJlK1uq8n5pU2a3eb5PXUZdrfqjQEDXgDmlJc
JQCMGw2yN/eop8XkHO7VTjSQSRSnhu515f+V7oDltzHthtKSND3y/VCn5W4OE6Ji7ysq5OQmd2Xp
Vu8HxmoKHvBy3rCO7jgEYVxSZJC/QIfwyHhy6kZpzUGgNnln89L2Di68knjhvtb7ajS4s47kLF+1
KU6Bq6penBubylmLMWKMImSe9grOBQjXVoRK94+Bh1nvXRNWI7c+TBAV/SE/SjO8USnt2atZIJhr
CFh1pPEx2AT8vNgsajEjViGNH0/c7NQz9YuWW5upWr+GjqUJ7TtbiNjZ+yWl3z+vUY21C3UchbV9
ribGsBk4iBSTQZNrXhmdAS2OUToKMzO8RWXkTdupmOKGfi2PqMHHdS8au2LPKqc13l2x6iyEP93l
hqRwJc8h2TwPyrLm6lgfkahRd12I3nXQka5zMf4hUddbhVlvn3oGu539lAkSpzpCHrTSGZQD17mk
B8a03GHw9OI+/wFJH8sJlNmfFMNXqNcHxkVA3FTGsKtV5xRUQhs23HlUaFUY7Obt+Am78EAgQA9y
LiO1Im1HBuUzIR8+j2Q/OmgzzCcZLVSDzcZFWwhv57cLA6dmjEP1+ns3QQNK51FvYBjyvqG9FEIu
vq72yehDTT90xy24Ml/4PxY2TLC/SDPHxRQ3nRFwpNDsLxrJAjA0inE4fjtUj8xY+pH0HI3KmiOl
T28/4453AN+KVUkUuXbes1Mt8+86BG+WibSlZf+Cm5xBIznAeHt5O9xRN//1qvrvDS5lHRTbjgWX
quSDvSZznAFP7+tdWZsNywsFoN+Qg67d+RssaheF6SMu/SulnsHnczJskz5ehsCfTN8GPPr9tCtM
+E+kT0oXcnDT6HrUPI2vgE3J/VAywUROHmR0eoSjsUcDpfB9Sfasi8+CbSs/HBi4PEfv4XyKQqe7
AbO4YoqWsc7bM5si9LnGnE2srKA2ltnu0zzQrAKEXUnNIooiUlz29elEaZhrv90vUWE60R0/m2kP
OexWQDn0V+LJ9c1er+9/iLa8zhn4KxByaRRjH8+TgvhF2Of4tn4+pTTy5kjO9+nBSmsoaaL6CQo7
5hH47RzR78Wep6Yt0qcj7YKvlaIWfaqYOUHhY47bRsXcniH4HCF2hJjPHVeNyjpj141xAepT2v9j
xIEGNoV67BhSxBqxd7nxqRYAnSzPBEEEDpg2JzEE0zvx27lIR78/o+UkfMWp+TukmCIEfd/tZ1mr
JhfmOaDNZXIxFhRD53Gahd5iUI3Q1m6pmsmbRwIxvq17ZPxhPQ4Fkbn+zrdWbvdCAZlZmc2mbuHr
LflFJRVxz+Uy28q65JbOKO4AFHb1PBG+KnByGITwZxIR+RY7v3LzHDcX+aoUhQhmfhp9hPoA4SE7
ALm/ttdrx8TCrCqg6fT23ZrYYP7DOuGtYYgE5aNsrE4LJklXKY+n+3JVwhLkYXAVhlIFIN0gUK5s
rwBmvcRvfAQuBSoQt+LNzZ5HLISXdJAZsMq35Lacitcd/ZrUL5jBJpiLYhtludz8M0Z0C3yFLRmb
GRrpBcqIDShLHPQ8vj4wD5PY/yG2/iU5fHnrTEFrszGg5GhIGeHAFkj3wZluEivAWX0crHOFoiWU
q1NTgyhUzehEptby4CBilZAJX2Xsu+YDM1etb0QsV+Ssu4PpyDSu1EP16bJikPhBw90CUhdmY5vX
SPkpDq6UyP1PEajQCjB9+QrbVApbnLzXrg1a22yWQA9uQTJcHDwzEM0fGMky8uw5jZNzpqrNXcDN
sl4/H28I/xBuo4hUh7G5SX33Kk5E/lR0Du1kJEhffbzVBT8caQn+jITZVEt37JKYQdr4bcmaP9Fo
AUxlOBukUSsR26ttkGi0jMb5t3Sq+6OY18Mketn/tuIUyXpnzc3YspGQecwyWzSJPWCOqLmwsRWZ
589n2iPmfL8YY9r1RqVHWdwrjr6el2CNKz+qrmDB6QGxRHSlTpPKvtoycVzSpc50rnjIbe0N4z3G
uUup41JqyUNZCPqhenFUiW5o9xVg1F9dTb+pBpi8PbcjVMNQK6gpHLr3HzjMOormc3AiFJvCppU4
l0j4DLbRAiT2qaMYHoUs6q6yWED3b4xYrO/8oKcVb328bOIDSTbkb5G6J8aBQXFWK2qKkr0nez1B
9eU65xZiHHpSiPC4bhpjY3h2yezaADhV7wCVdcJzQqU7JH0UHiuF73eDgDgbOxSkhx47Cqiz5G9e
iXx/lubwRr/I7HN3Yd+M8OveJUe0o4LkRW1wvC6Ig90rOSMr5m3WVOu5zYDPf71ZQcCqjJh2n9g5
tckLiZ5DCet0cLXovgItGArkhglLCDtTPWAp1lizixXuDaCZPe4FRJMZ1DIweuWlG8h4U6Mp+5p6
xhBlJJH+FOdZ5zIbridnU91uFJuviXSKEi+QJuolxcpww8u/b7CT8cASRKOdwd/oFOZGeE67ahnH
RgRudeSWuGdIuRP1xjBQur+Nz1SrO1asCevbYpMze9ctCx/aPH6U6PSOnbgrY3GzUTFMWTsCHedF
RvRL+9ImarTivXj7S2ibeXPen3kfecIavknpKFHudYcEtxtaIJt37fbwgfUtPc8/DnKYNJgqGVv+
xgW3KVjLcaOoNc8NM7cL74vHBCCH9wJEaC/f7Hyv1jk3cxldkcmCRl5sZoqrQROwH8ZHMZYs6FOa
gNQyAfAA3qK5475yQt3d8aksMP2vjtOW2Vd69QGIORcfk9c7k92Y6NIKZxv5oCCBoMh/rIFB4hWm
fHasJPZElqUDtIahyHNPAcGy7BKO1rQ3SDVRt0x99A6rjn6DS6FQ1BVqgGiPgkmV4GDKpHslANmy
V8UwGYlrUfiBgnGGkWphWk8eFiBCLLzX+UyIgQ09qUjDwWPRTAnERtQ5UBhRaqG7CsaWWns7vZdT
hY5091ptnxx7Fx6+7gKwx/SZDgL4aPEGM8gx8rZXikM3pG6P8jGz4M29rET2eMDuRRpCGOdgVSDc
RKJwBFkk/5xQ/Lo/RvUw7zdw5g2M0bpNwW0e8P9uH9tRKbhHttA9Md0gfAtGPDI1ZIyWOWVrlzUC
/yK/P5jxZqF1UlC11S9drZ/n64t8w9TwxAnmnglnowiO9ubDJGsnP++gA45rAhdZ4Naldtr4Av4v
UXlUhyWyCm8jIwjO+lg+t8fELCVZtvynkMcD+xaOl6nPLNl6jnv9wzECiO12JNnuASysSg7Q/GQB
1FcMtHyLIfG10UKnPSo6TQvRsIvDSCMlLlUNtByxoTJToHPKPnstUVhj9BuYu6fquaMv7hdk1B3i
p8dqlIFCn02iRt+1A2hqE0XJ/zdQe7fW0pDAPfI/v5yK4JF2ZYxXfvQqAu9RMgItPseyFfl+jx+R
hscVBfVo1tlsvae60jt01uGRE3kBDmHlEcHV14F5TPPMMqt1lhRy0FzAHpw/UyyA7L7wAbABe69u
tWr4pYFlIWDyyYur1aYco6Wt09FCyo6cmKSb/O+d2ygnNZx0A/RDHGBVvMUmcp1Vlfoqy0kk5ndy
VcMYgpTTQpRhiBVAaDSO9MS1KYQrPkkZui0+b0zbCyjJG93eaZDoLc5Eqfdn9/zFTpqUIMJJC0mk
w1uumLB6HzDGEcIW5jMU3XMSJLs8quT4AWQjZSqDc4LclhzYhxtLVDYRgBJLkBoFM6Znq505eG71
3310ZDKlkZjIdBIia9BaCH9kQw3mHmxr+EfUEgFx/RIVl8MdV/r7h8geWQjIMLXUw9jFa+FqK99+
prReuQwGrZrB2aPHl92L/QFWGuzbwY44cnP1tiveruFcGJ31F42KQNOlBrT3l6PmHRGB4r9K3tQx
C995opEn0ToEo4h/2iSP87f7vgjwMqHzp3220y9oDIZr4j9oxqHWYvIoTVOA1wiSy9gJBT3B+shz
klde1nbp/hPIsgbSQwEF5UBdE4VUajwvYMZa5mHn8gWJ4Zk0ys7KNRv1Yjick27iWAjDmZ+xtWHL
szWrexSh5f+aX/5mSF0FFyKqxshHgJhEKEsCgboSUhooFcrU9gyqYyIlu5RqWvfb1fAJiRhS+b2U
wlkSIkezhjzedPCjEVW3xRbtZ+GoHkns7rsX2Wn6yy8KLTOfarU8W21GDU7+r3Ncysb7ac7Jwr6W
jlQwMYgfyuxxTWRDy2jfbIKUDTooE2yskcseAWHRvOF45oWmKYbAepQsdnfDEwzc3i0dpr1wgaGF
/1Keu1OctMXzqpKnBTcoSAiQA/Ps5+8lGvwnGp+onzXcHS7IsSvEqqueqCbYVa1uuppSnOTsZiHH
A6NxfawsarzadBfVi63IBK5bsnfWRu1lXWqz+UDJaIxJuwrzJ73M+pmm3fVsb16ADcCrQRa2pX8a
NuRHBIqMVVL3b9GXOh5gWsExNoxBITAC6oBNv2BBFiGekUVzCidr4Cs2zIRZUzoDRX7jYQq6zn4p
6zfkfYfTIiOAOpn6FPSOsR8YEMG3qbm34DNoEipQFiPx9L+rsOgA1TcP0LXXwbpEmsOlJeI6bpBG
4S5ECYgV+cwWVRN7yOkrscbFCkjtFnR7HpYvyBGzbBcdTf7W+rxLJHngFohVlbCo58j9CnAi9I00
vCz9ikfLV7h0oCwQvuUz0LpMbKhgYBiLvSI/yN61gVIUDl+i13beny5sM9PNEXA59Leg2z+ka7ic
oT0FOx56bvBFNGJIRk2Tkg/2rl8S0sz+t3zDL0/eHO6D7FuNowU2HzxCC9b5HTQY2t7wM+HRT2m0
NYmD49tMuLH9u5ujR2OAxJhqkPX6DKh5iZbjecdL5GSbhx9xOaq4jOxgM1Yv+q8k2OavGezp8Btp
zHQaNGvNFHcp7Mi1T9p9ZSm3eRgM74c8MWbplYQZdaAaraeQ4WZ4Cx2EWb6FIJNL7F9Smc/F3WHy
PStKs4R68glNCs4WYH0uAjRx1OvzhhPmDUx1X0+rpGJrKxpq28RPbiu09qKLSGXPHmkTT+xEfxmF
LH2Bn1uSSd0XiofDODk3kJkF4hhu48jsOYB2iZvmIw9BXf19bhTiIjwIVPxmkNj8qAh2cVNuf5Xs
iIrF9icZ+jvJO3wH+z/slfwLj4l3ZXW1GlijP8J1hroNyydi4GJEk7EXJV0TgWY2iSLUpIwB9+6V
lr4YCvfKbqD4E+g2vBbVwwOcTYEgim1uQBQK/nhpWzGJgF1uTuVuxAL5uv3XsVEajO9QyXdX0eSJ
4HZLZAo9VRQockzjsCMmQkG8BhiyAAQos475t4w6jn55wIAdvlWJIctgaMgkdfBQWNS1k96me3+/
5eKuCRacTsQgJyNrVewUTWGdpfUoOh7EkENmMYU4tfrb203GgQfNbTLlu6E5oFW6j25+hZ8QN4RI
T9df4NpdK5cfORv6mHTnCTIx80EqV0H4n/A3FBXgBiq6wM5I19Tw4Z9ul72F+U5OJDDPSJ/idM4E
Vy4PKEdoSaLCjtQ894zXLLKybbIjHN770W91MIfCKib+E5Me1x8P1nBAjuqE2DLNJWj+/meGJUz8
zFzFIDg9FKwlfYV/glU8r4EUgHrLqVZKx7HO4Vsh0I8ZP9VaniqeVDcVH64HVEF9AYmDHq+NPCAw
OpmQjn+5u2QBQM07l7D+3Vr/c+PpcuZLZwhpwQOvDaZ6OBVE7vIKjVm6HHyyOpNOX2iKwW790LOe
+XAhjoMN5NGS1/vCMpZMKh6UV4HhNIVAwpj5sw6v+Pns+/zYtAUxavWjKTulnDJZmrAQ6o0H8n2i
WJz9g+Lrp9fQLJCRtT7vmsYyXAkAZz6UCEF/NNIRlW6p9nE08cBuLz6x0i0NGvuNf+U4d3oXkh5C
S9GZwsviXhfjQfcGQangB80Aggemya7/8w2MUXKgFbjeinN+1CG//mXmoVmdzR+SQ+cKhkIzDguz
YbSQFBPzVBfmtdmQ7pN8W27LKmOk6X63THVvi1YIeWYxyFrCivyfzZHBKzP+kKuvYvIJSY726gqw
TuWnwcSms8DPQp33whIjO6gZRv+0ZN+dpTHuPGFUXgZ4dUlBzlcpZmIjZlvezP2P2uqCdZghPxXO
zE9mP9vGxmRTUcR+9l6hBw8FOAF21i+lo63hA0vdahIL1n5tEuWF7D+yKcS+INh0vcLlIjFTcjk+
O+4c3DeXMPIAvMipld7pipaD5Ez0Ey3wkRHu3QaVypIe2OueTLn5kVCKFhZ/9bPoWU71gxalqq9j
DnnCAD1MOTwZTBZdvvFbknwByLILzlwOfsCnuJK6XIDe9JJL5FdJEKi/FqfCSXfrALKG2uzCfxRf
xIkerM/xaN7mHtw62ucNe9s/+FGrrz6CxuC9OSx/PeQbAGW5IW2N2OZOTroY/4dRd2amc4tWQgJ/
NvwnRPoGcEiGUtYJ1nDfBjpOLnKP63RxgCC1lcNd4R3zu48Zt68nF/8j1+51t/1Y6AtDOaXmeJFY
2WBZb6unjJFtnKxuvU491q7FzEL62l5yAJuUckfFv6qez0UB6AKETe1ZYuAj+3ubOvSvSLgzrZZs
ceucbLcXVlbKLmnUOvTx1cv/2JBoy7c8RQ5FwjEmqj+SJoksZenbYOH/hXNlgbrIYOq+5AG1nypI
YmzcvDelqOS/WqcX0+AiZthGdbo+aD05+y+T2cz6Ge/LWlnXxUxwJJNzUrN9Iy/Bkx+RJ1IcxfH+
MO/D3XiVzd26eSDDi1iFXH2Lw3+UCrWznal3RH1kgJrM89mDDNkrUr+a9R1zKo/A9XYuD8qgBQ1b
3UmhQWTAT4hLx2xv9Bdjuxbw2a9PVXzY1m3yJzCDneXMtJzImdqOBj28yMTJ4ETekSk7jJr/5xXU
pq4P/YYODGZhUYUk/oepQAkxPh71g4OUTT03jzHzat5kGVU64FK7n2F9BiSZddoQ6DDop/rwKwgS
xKbqeP9b4zfHNtBWlDoUmdvxaFm1BCsUz893dkFj+iv0lw4Q+tn9gdItcSJRX5EVnyLYAVbbMSss
ngaZBxKW0XulH3MMfg3mRDC0o+YRYASkJoSOoHnDAkpm74NcI8cCL5quJAcqDtHQ5GnYyFwciEju
Mm+lScxDGltmaPTGyavyxe0pGp6HZpH1loGnHP+97/OOSChhmRanxcP21Bx61ZBLxswvW8Cz+phR
Itu+wECmOim7Xsr7S8ns052L9aNJCX01WPJ/Vlo7UG0Q6CB/AgruLpN4LmLLLt94CfEVJ21Vk7Fa
gZCQNW8KxyePuY3GwXpE8ApUpy3YMjqWBtSbJ9KPEMd5KGADqSQ3AKu9UYNpfh37xrH8kKCCBK3A
mpKFRsQ2KHqR2HOKpfNvdE9+udNw2aglHpDNDFKPmbz8KJiEih5XKLmY3NsAx3Q+BmhUflvWtKnR
bH3mgy6tFErl0SP0LJGnNLmWLz84GfgT4n2u8rgTZG28Hwn434i9VDg5nl6oNHZtZQ2Pa575vHSX
+mFgQSRFtYexXEHNv91JssFvo+ceo32OZkTiXiwxdQ+sBhzymorXBYp9Ed4BKtYPx9BJJ1jFzm5P
aFyAkxMn/BpAkOC4qgYLkRR72hBZYRzdIcncPaAE58kVrd2Vjw2zBZu9H43yw+hC2slwfV+DMNYI
/q3XilO8ei+StUIglq44r6XvN4ixwFdtlneM6FX3ChM06A+hGwrREv/uv+dcFozh1h9p49tltT1U
iTIc3LKEdi5j7jYGLuMdxoR0mNJKqiCJgwugrGrjcryJh8coHnbGiias6Ixxq/kU1uwYUsQBsrUA
KDMVBrbGZrtLcaLVYpzK4I6nInWhjgmxvAx7u/sxGjIauRS8Erb6YW0Cs94RZ5jvf6GSGlfonqLf
4QSCFbQHXia970p3K1XDcxdVDAx6PRIlg/cpmvuu5C0dc+TZLHTd3stdfr6T8tQ7dc4/0ZFSm28/
+peSezt+qlSGkc2me1bWJp3JVUtrTVtaSL6s5JLYOMrsCsZ+dcE4bvOKvGs9DvRzvVxpH2rDsXnW
JU0pqAQC4K5PgTG7bS8vb7EywFaJfszjkWgVcUY9KHO8ddB3/tqTYAwXfPHvlYSSaUBYvRfL8+mV
aj8ECd94w8oMLYh6L0SCLgjs17WvB4ShrBbfGDgNE+e+/i361tbgMtSHvToRy+dWZ0ZzTmVn5XJR
+T1xuMarFD9T5bynLwfi0AzBZASPdvy2tHYhzQYx+Ks+TAehLmbaxWian9m9jJo/8j/ihLgjwtOE
Gp17p3qUWRbd2v6DSS4YD89hfabnWIodIoHh4JfKPYJZO6hSaoyUJCGQGQ6brwsohVtTmMerPesn
e4fV4TF6RDMFK9kVO02dtig/cNASU7zU1J1Kmb5bZLkOyFXADHPpzufB1gTwREBLmLW3CTG9hpM3
ZJGPG03afposHnYOl1yhad/c250mbiFHfoFUxyBDryON7n73lpMfyvA7Y7hs4QATdBLy5nM9WgjF
vuFpRxCnEP7W97LTq6Ob76Ig+zvkHZCT/W+dlEFLi9kViev+b2B9HV55P7YX0Cl0EUExIlb1kNsi
dSbreoYm/rFpEvo+ZhaxzKb7DDgCEz+TnjGLSwuZjGLBImk6MSD9mlxZyaAbWO78ogRgGfv14LXE
lgLF0NPlC5xhfbMv4qb9CznPNryWdBZSuOYRUKr7iXbnrIPi80yOC3K4a9jcFNIh9I7/wmM7HA0A
/1JKJg0dRQoCa3C7uz4xEVJ7sy05zdFyw/2/3Hgl8MfT09e/uTKRS3QoDdOOJRnn31S5i3Zv0YmM
23AS0SwQPNbUaupd7X2SfdixN/Lwpla6jEgsRfhPEJqTEyUHJrbiATVs9TwCskpUeKBWm/pmu0PJ
XsI/elpGRbmbqU19eLSoTLWUHiRr57bbGgUbJjjDz1HKWq53pgK09lgL+0CcR6eq/xb6pVHwFrib
i7wiRL45i34fGy8nTpYVesXD2rY6JAJWcoWlJOdw+TyWbIzRrNiGRpcC2qcq4F1bdfbJmArMX0YO
l8F2uYNt87z9jnFFzIJzLON/A+VmAJGMVkNPnrXyZ8glMaPLpubfgYXu4xyzpM1SGBo7UfRtG2e8
2xZMU6bQ00OPyxxriDCJat/EgnBkWsGIqcJXHp6lyq+NF49LldF5wWKxZ57gQsx9S0QKGwUO00ql
XI1xSvOZWjjZRPeXpKKSi7mmNcK42hMFRARNckq0VP8qRl/Q05S4Jd/8UuLHk8NJL/w6/+fHlUkG
BxEYV2TBGdg5662BvGNkN27UuasVH7QH7OS+TA2II8CpFlgmLqa/F4h/99c/hkiMrY+zhCLMW1eY
RCHKXaMbIh4lBTO/FsIQZYkohw4249/3oNFRR4URvQoTht8ZLmIvv4S446wdKwFTlQ/g5iPajFwN
BUDMWRl3Wq9ZwneFfxskGdiSnQQvKvQdQfi5GksH0VO2qecKufOLY/VxAFpIGBZfKrYyOdAuJodz
z+icij2nFADzT/3vR2PRYxboADFVLP1pbzMcDh4WHSInykxykBBfpirm4sEJD2aoHlG24UdG6v7o
JbGl8qVOHvCpzDI0MlZBJCqOWEyjYn9AvrkalQiIIakxRG4GVU2NqREgAaCaE1DY6er05qsqKqEG
sFxXh+kOFPxiRZyb/jSz4Y1qXC+0l8zylVhyhrNkwBYq73dF44siNhvsOvrIyZzG7OtwILM04lwo
7zMMivHFhA4tWQJiYKyGNPMtZa92tsescRGexqzPn2VT85+mnN3I+HsoXivDt9bCw9U2mfbKur4t
MVr7xbKfOF1FhSsTxGNNm+DJp5GipAVppJFxkmsgS9tQuGvM8beVfnn6rm5qIYcEhkJOthKir6AO
8FgICwYkJC7EqGekLRWOg9tDDcuXTfh74Pp/RU10rwRX78vLkcBzTGruHoACPcvWPqhMAZZLHK2X
MNBSW8H14922WjJTL/sJR+UIEDunl9EC87Hu0pUOZ8MkfG1IGmbqP5mDHcTgVBeWWy+qSJV+S9ba
f+M0aym/Lzc6eLKQ4U9b6jJllcuKkBN8z/9ACS4KkFiy0/UsY4B+MYpR2abU1W4VSxjhFo4P2+Wo
b6o5aGiFkT56W/ASR2N+Hs4oD0QeZSQQExlSE25aLIrSeW5HdIKBiOivO6888QmNdxW3/JlJOcq7
MsnAeJIWjGagzoeHq44B0seujp0XvwHFQ9RqeCeOfXpbLRWDod6ez7Z4MwkjL3Ha4FrXO8nUAT+V
O4a1EHyvtp/TFwPxMFEdEOVqFl1NT+3HnFlq3WRh0yCi0d52r35htdode+Q2lRCyBiM4ihug4b53
seeFcgXsVoOjiT+Q3PS0ExHVChKGaxuLW5egEV0WOSqLs12Sv0MMgn1/lOq83/Yt/a8GPXJcwLEI
ILFQ8MDMWnk0Zl5MYPtn8yNNsK9de6c1FPqTJ6b8GHHG+06tk1wittB9oZO9BKVI7EqzToOOmFRg
lOm3b/jZyDq4o90uC18luOWCiqlLlvcesvXNxIYLag4oKTb0WMhG1oh+1Bd7kC+YG3akXIfj9Bp1
HaKH1XZlegYt7ENU9nGRybVX+Vt6UrHDdIF8N0f7+7vrE/Y0oBaeyQA6JU3fF66dg1Ge+va4kMwR
wYA0MkV7Jsk7jTJgIpFos2oJbfNcD6xqKUra3uLx0YLjA+XEDNIkMC9Bsmd2tFCqMCnt7Z3gm377
GB6KrzJwWqpw2PtBXWRIsUC7UjoMn+QZNnZNzjYio9mrp2TDT6u8RyXDbhW4+9DydqiOeKYiqtbT
kjoIy6fzd7QJ6lM/etyYXvoJOmW/45zjejBnzz0PCpDKOaqboSGCMfV6tV+j6hc/JzvvhsizOkAf
SrU7D6Cuw/9jsEORk2/1kjUpOfY7IEee4Uhk7mMq39dlohdQlCNvfJMfV4P6m5k3FPBKuOhCBTKg
36h79XbNjeg4DymnbFba57RmWKXJUmZgZWl2HuiKwCAGer5EQRid2426vll9s99rIx7A0BRDxuQA
dd06eQtCaoZhr52vC7VW8Qq9E0eMbiCIlK0+ocRs9NRLWIbp26iMq63a4x9KsS0BlsECV7VDGq1n
WpOPOrJvFX8X3zemY48YZ/C3DH+yUXNLncQUr29Agkw+ax3VASWvnv7dE55irF/PV158et/kjYfd
61RMxmFqOBpoMM/wap4kBpXBap9aLW5HWpxem3Nv0f/grPWP+yAIZtnRCfNvGZD3k6lnewdTryEk
1c0vphy6EGRfk0oV1jaVOw1lpyF+Vr9Gq6KWONkXpj53WQNh6JzznNThycG/K40s3uWneBgVlxIl
nWUXzpo4wVr/tJbm88IAWlkMGy1NLWG2iyVm5Aers6m1OkIEP4OY/0nIJWtO4zKSTWsJtr2aNKiv
s/aIwgNAfE605KTYjGixuq9lglM6BgzDm6SFJ+CytlLoodZbZKAAlUN16FB24H1UfiZhuTi7gSCv
8PDMUvfAiRCMrY+foTM6BkalUX3eocAmp/2G0JfRuueiWp42BjTqQvHOsaLsWV1HxuPufFQ+bJnT
kCLDRYKC2njvyNiG7ksbFPPQbmlCJD5xDcJApfLciO2uGWTXrSZuRD4Bv7bK26NQzg2noAn1+0ax
xCsTb2hTSMSYa9RHlRFKTXDO9Xsb0lA/Z/j3x3U3EtjBopaNBDOz6rYoWKT6jVrVqfv62z6PDDQz
/Nu+5VExZ8/KR2pSaGxuOi6WBZJTTbTnlicpQPr0PRu92PZBsdYCLFxOhETmZFdjTwCZXDHs6Fh3
21v/hSfG4y7ej6CGeQjSZv8MNt02qx2ZByqnpYxUKwuVanRZBtarjlK8clIlPH98xgAYpMJLERPU
V5Ao+YepG6zLOzQCtk3iNQZRFb4RLv3vj05fwPMck9p+owJW3qiHrQwRVNe0cov3wvBOZW3yZVDF
UGgou1nH6JsnGA/Tt+3X4fWP/63ZiC8xza6Q9lPxguz9Azbkf3mke0kAQuUb6VsQYiDsMv4dk1jN
7pPgUjSSMd25b9D/siI2zmn18ipaeR4AhH0H02wVU3BW9j5eSk7sk5v1C4RIYx9g4i61vYC0a9z9
nzXSfzLysNO9vqpaPUQlzH/gcewLJxnEky+2nPncH9EXeb87F51Ik3ykLnoypMBfM6xFmBy9Ri+C
2tUWDWMdgyx8L3Ik6mpP3W42ihXK+tjP9nocqwggIDnfPwbqibnYvwqIb70uT2j/3TWwuayo9ubN
7kzhJoUeXml9BnC/JnwIWRGn6Q725daMvsch4zGvlgJAY9MvpMwNpy72Kb18OpkFFjiwP6lIyBRJ
KGWvBNDt7848EFK03R6x7UIuRuulMimV/S7bv8HvJyY/I0GGHG8mxP4t2TTS72XQYE/EdXCZlSfo
RDUhUsRQ35SThfNPg87cfzD5WJp4cEtonOqYoXP1oTQLc4G3b+4q3Bq3mCIPvcjWnkrZ9927/wDD
8YAasbI+5pzBD/UVCO1ddctcH9e4DXAYFU4FOl8xXJhda//ebWEBu9/2oVXL22+5gLKdpF1M+Mc5
440APR8ALP+ufnS5PyvbyQ4EjgAJ2apaR0DRmt2Av5ZGAp3GtPFpm5pruYzEynOeZqehQKgoFW7C
WSatwkfJ3DICp+6vsedhyz8sEHgqn4Ydb+oYJir+v3LsmMnp1/WOJFYLrEhGusArif6wXFuW5pGd
PP0I9bYt9WM4iTxc1koIJYqxzm4b5iW8SpCiCrYb7dyVEZmsGWzkVw9Yo8CJRU5LHp76+I6mDdtc
DEUNcgEqFchK5eexNVgY1GwoKkqhTBEYzHurpy419mSyeV1N1a2KoCsPEhbGkgNF4/Gk34/XTBEF
l43URAI8W3lX8maSEe9NFcbn6wolWg6Ff4I+XBvafbI3Ek2+5C1XL0gRk2uf1ppeaUAvZPshUotT
Exv3P3STBVtDa1ROkgQV7zHbx4lEUkXzNGGvP4g89P6W4BR3g5w6Lvzdrep5dqnVPgrcsHoOkmfP
2fdTLtlCgHFauD19bb6USY7dash7m0VHYO13V2WvCmm/JQLtI1nfu2FCkBNHE2WynTKpbENcW7f8
7uzLj6VzyAdtrrs4jPzC3QbfYC8PvnpijBjSIpZ798i1yrfSNJHiwSQ8oWpgbZSvPAN2I2nHruRg
tzmWj/GwbVaviUNRVFmPMQr6FulxpIxmGaC5r3fu80kHSjfFK8DSRPgDvwuyuYJaRodTdB8eTj8r
uvRnRMv1+a/NeHvCdgmvbHu1LzyIdQpe0sw8gNWICFqsO5wVRI5Fk5xCOFpb+R/h//RFFvkwKW4J
6pY4lXGKvThQtybtbsoGaE+IqTc+vkwsh1oZhSc0DoaYl7KUsYkyS7eBLntERAl6j2DbBG7QCnkO
z51AvcQRnz5nDUePTYe71q5BW+Y1rj4fN3/UU6HV9XGU7PsrOYLh9QG3bQTb+VuyKMU132tflm4G
GM43SQvGz12YWLvsfMVmm7Hc87kaX6kWa5obS61F7oserVv52FbghZiuvXW1jjjICFeIPPQyd6DU
CYschsY8TvCQdB6/LXyNlEQM0qXVl1ATdT7m1+LvkF4zs3JqutHGFRVxaillcyGUbs9rH8i2fJQw
K81dL8RNj065uJkQ3k5zgVuMEBL1lOdJAUr/lP6YVRAub/oFZRh8lDh4TkQ9edaLFBL+0Akll3Sl
EOaEjFShhJoajnKU1F38e6LhfabLiqYrHOL1aLhN6PTr1M5mL/GRWcrrtCOdXk3Xu4kvfu+maMQU
QZEj7PpoOBhT0tXvWijQ9yPVPCULp0aWa9oVKfjb0gYKNCSPNy+l7WZJT/MTSa+SBFdcJepz7W2Q
fXC51xv7b5KsxCv42Zyy5vkgUrKTXkYkH9TeQf5YmOtCytxqVYkZlQ6Nm/CDk2lXOjfSlEbyBTa5
YefNZFpqSG/7haZBubdArXn0oMPLhGkEgJsjoY6RueK8f5uDi1po/IDgjj/0VqgCIgzF49OiGiT8
mm6WUKbVM65M+ZMz5s7id8Vr7SqriwLLmx30EJVLE9m46NTOVi63L6g4TBdut3k9k+U4njyAmHts
vBD29xon1hu+AzidHG1uPxnqmMeu4AgA10cGetsnd/sm7OIGtmeVXT1AMNuqHIOCOJ2jcX/5aR8U
P+L4nA8rK3TNAwzTVg1L8S2+3SyY4SDoXZaiAj4c82Sc8m4KHIBluiPCml9zdsiHY2oY+uWu2BTN
KKzki3TJ0+vEQP4E8QjzeaWHPfikoXBdn3THNM3tS2qCM+nI7qU4JbABY6Fm5INh1pXKZOAf1kkL
CVfnf3ymWy2LSV+KPBd7DjUWA9ne/MBhXyry9C/32YWXQxANuP6C5F11l6JnXcLRocBzqT9kaT3B
GzXnEboVN3U4OSihoKVqSheQpSSgb4GItu/qF4u6HsIT+oMN6rszuzPP2pqFhZxGCak8VdoXoKfy
asjjrxETdMNes01TYAjUPJGro20wN2QaM/c4oQogQCqqLjVFV6OgDaShqk57+HCHdyoLM+umcAax
wD0Es0p3x1Lsi2qqV+JXBhdjwOf/d2XXEN82nMxgIwM/7PmpvzPyUh70+3Je0rCT/e/8UBZskOiB
Ig8IItuQuobazYgpT2Gdqr6OiNEE0NK9kdrEjO+E7/rbpVNjcxe0Z4VuE/R96mIi1NpOeiqtyWjJ
ALioPnJxD2Zkc2/0qTs7aowv2QmO21wIuyz8SK7Sq8PSFBN3RsWbAStbW2AKVh92n0t917z/5hER
+hivGJMyfU6Yd1L/arJcfhxG6GhB+kKLwNPqxCEKeMSN8qcJt/irLVLYtllJS46mET9TXJsjVbAk
FGJ8pQdQ3XpajAn8BooGwatbIygFnDoW039PiL24yKcmYs6HafmC5Y903mYNzBXi529LD1Xjbjjl
vQ8M8QSGt/DU+6vLQPZGhTGWSCfF9WXqacJg0IxryLg05ows/K2tFTs4vgoVVVBNCzbmf/oZF7TS
sdT05LzQajOTyiW7sy6S96qEGhXiS2l83gGdzB5iv3WjwMttsxeuVlSjOEXpMCE4w3YwpLbXWdRD
UeYTNooNlEe+5wE5oKsjVJsTZMPUYFWwgBtCfHzTgUlPl5dCGELMHpm+dammaRISHnzwFKKAjZ9L
TgNNJgcDnYwnIjXPtYd0eJpwaFpyy4rKCcli57oYq9KoBLKIZpQuCtfzoJv6vx5Js6g2dFkHCXNu
s9/CLTLJR55feP1L2QohBxxPUxRRBd5Rgis0LDMJQM3FnL091mJeFmE5XDspf/ILa2UZX4VP7Nsq
iUeFxJ2FW1rA6v0TVypng8fctRdOU3oTiLKD7fzmS88EQ0ek1WYQ/t7EPcbFtanja7rV2ZWENXN+
k3Eu0W3war6+PTg9FWD+X2IYB9cQG0WFYMl8Tvl+Jgwcr34wm8T3XalXSfWvGMxlsUVzILDlwv0y
Y/WrnAPlv4pblD/CwoxDtGhNXoGa9BybRcfNyDbFxJQB1YSISJojHUgesCbAAnWLmjjjhXUDbp3B
9vBL6+SZa4IeOXNKMksSS01EH1adep/HIne7N1WYMqde21aZc7hUDW0Lq0aCxRbEWKTv+hMempS9
Au0IPrmEQHTUAYpnIzLAinjI6JLwWd8J+n0b6x/bAND+PPfxiQ/6sF6wagi25E4djWbZGEadAynP
Ara6h3RlKPfkpBXw3ctfGMCxX1JCE/PJ0RvD2bdhBz2KCaeKRcHeb4CsxkygV+r7gGoXHKh7//lJ
mhp9Gre9UOHGD3TG7QQ5IlLZi8YkXfDVfs143u5HdICey2a9HaxXAfD0Ya1ryZSUoPBRos0vJ2mC
GFTSgKAKdr/UzNgn4M3dyrogHWo7sEO/UfZjd3iCFzSHkK5p+d3ux/jwts3ZAjBpLg/4osi8WDcf
KwVWqa0VCP2Cb3DtLNZbF+DohaNTPteKyhkNA+ORYoCGgUBqGR2odEBYYWjXanO6sjC9/LbsC5lb
mdFiiFwV08svUFpsKLsHsZ3mRguh8asCXZYTKc052+nosuivEety+BUpz8/ZWJsRJKv/kkLLep43
7lLn6oImv+AIsyFtW2o63nc6UlRMbe/+p1KAUlLniNjLh3px8+4fFQVZ7di13FibeDAymQ+1DSZN
u9VptJVaMt3gmC/o4Gy4pUEbe+ytAM9xsZSlYKL1FAjgykujsaZ60r+Pud0fURsgP9O8GoAHddwe
mXw3wRRuVC3XfvJ3Gr8Dpcn3gJT5i+PxgTBJylyy5styB3rxBm9maSGHNu4+5zn3Gn4KjDHXGrf8
ndrgY3LChNDTf4ttznpW4QE4dm9kXuXbu7eFWBeOhThAbvOnT+u+yh0Mhl5fnCF9buyNVOS7Xa9P
2bzvtpI28qQfrCu3yNihFAnQCEKVmmBc+tt1xF1O+cVg2dPDbQ6RHD1rJdn5KTja+S9yhTDldcxp
LhkyLTzoPvm5tbav0lrMzpa3hC5U1sD/3CNHLAiIdzBdV5gZ2l35D7nFZlxs5URrmOAOK6vMMPHw
NjkHRfYfzxb6S47bfssETozmylpOPKDG+BygwpSc224UJxziwK7kbLosgoqY0Yb25MgI/PJo/Rrb
Mqx2Tugihxg0VJa+bA5hK55DJGuJ2H0Fn3kacPLhjVu8txRgJgtkCyQszwcUSVH32BVZjNk+96nw
BNKed+MgHoqCiZhTw3Qvf3lSw4Grb8Iw0arGDfyXkdTrBcqNhQJNsS+/i03uz8JcD4++qKqoniLF
NO4/59qnXYW/eQueDcDruxO60JP1pAtV4LNwyfKx5sbgimyS+B6QV/F5wD1BvrK9n5xIZFCoktuE
H3xlp/JOllEjt/BEST9myzaPmRtGfmwjw3VSEbHVR0SOAP9EoFKhlJdVEg+xrg+eXZOnlMzruSwo
z0BzlNw332SsHqg6VBvn21xnkCFtJoC2Ihw04nz7iUrhkHPjNjCgSiXegHpHVQrnYDzwdiSYqc7J
My5FsueJlGN43OjIqRTfO0YTYV2fI5rn0D+aX2f0xu6RdiWwvIlfGrNL2byRUZOssP3iUOll7qlI
oDoT2wVOCA3dnz06iLU8WUFw0NGQ7FvrSwdGkg7DuSfEaH6Rb6zAAYm7+AvDmwxUI/3+zCXkJtY/
k080ZRdQ5TCyJXhS9S6bLmAcc4hPKBmpirc91YFu7i0dSRQLqBwsGjjuYlnpfE0vVjJS+SYkNB9a
UIM4nIl5AHG/btPan4g1hZlpOmUvBOiERPdRmo7DhpMDqxz30edp2JiniIVDXkhdem0IMYMUN5v2
p5o3oq43H9ZJNJ7AHOEZYzamBnwWuvkNBs1g3nvk8MW6MwAADemLpywXb7JjAtixg49jp9NY0Mu8
Wiacy2DnFgS0UDJgv2tcYKXjDz/sOd1rmY/0m11lv5dX/VOZdlubs4cSbhRsvFtsS2w/Ea1HXQrh
jdrEwjoOu8z2A0zxZUkZ7i1NRO9VJnqn3xsdGkzG40IikZAXf1nTjct77XNssP4zGaSuDLbi+O8x
8Ky1cwooT9E4VDKqSE88iQv20phVnk4nha617ZsobWthM9I9L3y6r5UIgRsUDT0MXeTmMkE7RuBQ
AwVbuZBrwKU2WL7BPFKJHfuOl6l1yQ2m6ZtxkpVCNWjiIpH8rEGHxt4rBMU/AcG5UpUDq45J8oMK
v301cojJkyr/wdm58QFo8iU4XbbBfzF972Yyw9t2cMRZbdeIhJip5YzxPvPuqxvkmzG/8BwknDkq
DgVdjzTj770mmD48zjANfihBUw/jk1XuHmPNwzEVGm3S1otTllTaLuHed3N61VraqIaJbGZt/iuE
q86LWpch23yqK0g8apX+nmQxxvXEx0KNm7jv3pfYH3riocSEh25UqOsuGD465nVdfYB+FqgIaD34
TsX4WyaF/apPYrDjvtniFD/wkkS2zK0SIuHO5pHe7BDhBp8gCkOtoagtbUdaBwzfWPqgdjfMkRLd
Hk54OzhnW3/9QtFgBcPzTmQ3nyb4xLKPoVIC+HiaRgDzvJ1NCcu1AagQbh3DI2KTBqyVVVKDoUy3
uqgz+7IhAXgBuYV/NEkQoGI/yrxcr6aP99kQfE1OXG/vGSrTTSGp3YBryj1qUNroKoyulrUJYzP8
ci1kLPWWu0uWyS+nhKZWkHp2nhgRf/gyhN6bHN++vXQDma0ncoYzJA3FBUiCALuOQPGVDzaYADKj
VWWGVf9bVb4vfA2T0Zt4HcDaye1K+bD9gYmjM7pltFfMyM5C+1fy4ADB9hg1f7dXcNZto+VY+mAD
4IiQzQYk8ACZlQxU2BnwSZjflvrZ92WqKelFo+ZyYZGgGevJ7N8nqhATTDGvYvKjGSTar0cYtHjZ
7WEYvYunHyKSlqkFHfny3kCtMc2Vtr6TJ5gVgJ1gZVwKbrJJlpFKDWPZcTXdJzCkDs4PHNQfvmZH
295U+MiC0AK5LwI2E+7lgDaQc4X4KFvf84WcCJsJmkDthOEwzzIOi8oMc2SURL9t1bJG7iPKAd/0
NADJH1JTqKkb6cn9tu/BrEzCPuIulSnaTFTPHs+kbWn7/+D842C7RK3dyg0Nc/n0pz4CGoJIWhQ1
G6ci5KUDhKDRE6TEJB3vKOM41mARDh3BJ6aAv4SByfxpoSbq1+y+T3nathdJSTYeft95Hxe92mkH
cM4KKN/LCKbEvJZysu+yk6dNIxV/iMJqHYnigGqM/gxCIUTlJHRKkd/Dk/tiVqZ6hP++HjQMmeWz
lsA6z1I9eFU5qkpzVKSW8FE6zOOJLAR+hWOjB7aAntC9eGzcok4N/kiqYYugei0qClCbdWW3z1a2
YvESv1vKX3NBpxXY0sa1lehlUaF/OxlxWLmZ7WWdF8JE55XEcB78kF5UMEpbnk6n5Z5cOUuDajq0
fYjapASGDhM/0vNtWnr1EpLYR4N+FLdrs40QT3Rdebi2QLegyqow98k9ntdaYHWORbC1WCNj9WGu
PCyfwf85z3DTSPX7cYXZRwNN65dWC2LXKgPsC/GgCDV8YAU3JlznirUmbR8yNYVzOWAY+eKEMkTV
ezGjitB3qqWkF/3o4bCz/cRzxbWSHL3EjvadDAUe2scqZlcPURUw1bvvhlDEeB5GrznaK+svMrsb
Rv9NaskzeZO2bqwp5e6t4hM/a8JofmYnFhZjjFGYod94z6O4+39ULzascgdAw55MZRfRZ+EVZ7gX
GM+ME7Cnbkp8AnVwBQqRv6q3aI04oXJJBWLXiAtZ4qPVHBbs6wgONicvN++GmcyWbaeMxT3Nf/WO
7ozTctoIjsi0o61y/3lUKtP4JUR4jbFvrz7rpwuxswP/uU7pYeG+xfNor+2LcBe7oA70BwMtwGKD
ZJkpc1p+t1BymhQb8r9IS20zr5dohvyMqffCGrupeGptZs5gGJbT3l9IFLSPsZKJpQJq48UFfed7
HTABTHSeILVo2YAEeVs35hOXCXj8gZ73lSQPozx4u31d8ZEJqtQFKIHRrnhZc3j30SOs+mE4ZHNv
UaciCrN4ms0PqsCp73BUmOk4TkG6fIvhTVDjzmDiOQZOyIUDijIghWPuPkl74R/9FcTKO11XEdYR
6ri6qIAx+5ifEhw9fYZIVruk3m6CiijimChRC7VOh2yxBhLMd/AlOPm4N8yfYvNnJ+Aufy+KgP5J
gxH3ZDaP8jCei4YBhtUQDzDBBVA731d76y5co6f0IgdeaWMSmiIa81oa0fGpSJlJvbs6iGSaeAp0
dzInK16TEdAjojVSKK8IbNH6rDfcO8mRTMUZC2Cy3X2pdB5pjY+TlVmsXxjgE6XDZHmmxJFmmgJ6
/qROxt3zvIfbioCGZJB4D/zNayTuSTEB5XYXeY6pu2NmzQGw/oELpwDP98NN5I2anES1YMZd7XV9
ZnydmTM+qevsnlD/ypgE+WUWWw8pL0Oqa0qON8T3awxBvZ6ZwaCUagAQ/LnyiszDmU9+ckxvRPgp
fNNOS/Nk13Z1aX5QkydEmlmidJi/4+5XPl3pPLH5eWCyWqJwfe11cWLTf51f272UiYYGAefKP9dr
CgEyJwjFyupT9UVkoxqEuhN5uxqpSDEzvQWr9764LkiILYFPjkEz++w5JPOz6hX4hJPZbKvXYQl5
Y2LHDYRgf2jtMgb8iT7mqzlGF7zjxLDrDm1z7IY9E+dWLG/t2nHkqA/FuIXkrmiKcX3BZcze7Qsl
Rgv8SvoyJMg9ily6M0MB5lSH96yZT9EYBNF3SxSG/E+zLkhC0AeF7C/z7H7U4mKfylu9rgd1va4k
Ub6oSGUuww5e3a5m4KWWAeVf2FS/S3usu4VyV40u8MGXAv5qBRiQTdDioBVYS9N4530yQm3sH+H8
2lEo4VHl3sCkUaiDskTRFrjXa79LknDkY/u9kFMjUtPIbAbs/xqFfqh8nMiJMVvzFZWe5dg2G5du
qRmFZftHGvtOQ906scDTwj4iLR6b9zmvo8qlKYrWve7r8c/kNRY3a9OVmxHxITU+TGMmIjMufhmL
inrxOGb7P7V6q86nrL9XZOioASGcr0TCXIPdk+hgbjYv5fYue5bPvGaaPGgr7lNwVw1+1mu4n6/5
ESsqBqWrNGJnK7IsqdHC44mj8hmQf2reIUfCOGAHl1weLFN+q1yu7EdVutMgogXPK+uYyxOCek+R
TALsupfFCO8McF4kZuZ+03QKl3KOdh0J+j0inPgurEKQAPEGVXlzZDSrK9IME1URgZXGqgNUUXAa
OssU4v/z0v9szu5y5UGA1vHMI8RfTC2UNPZjy3br+DcKLLBXEGTeh8k6SZEZaEZa6B06rKh6/9iu
4muR9fr9+rJscj+7KMOtuq8ukbCXekgVd2BwHeO1WjCeCxXr9wPBdfC81i9F26qQIxeJJn6KChqL
SCQaq71ZC68lZgisw9N+/QIB0J9FxLzRjt2fQMNP2r3Jywb3YwrgHzs1GAyOrfPQMyk4vfExVrs7
VT9fDfHNWfG7fqevjsWHm1PRNdIu345KqWa7Cf7OHa++3roHhIiQXjyz1YsZk11VZqYEwaEQaWh3
yKuh4UiE1anNxsEYTuBTJGvHv9xqA9MvPHtYM+Th39hckwx82V56otSp1xsg9l7+p8K7H3TZVVnE
i7fYKBVmKI6AU/E23Zuh9XQj8CD3r3GDVpwg1u2LgSW2VNni84Kai4SYPhGqucAZ99goHA7XTvzm
FSrXAh8Y2u0EE5uAIwSZeb9/CboVRabqC3IRHF1THXcznzRG25AlFL+PlLWlgPpGzM9pQRwIMbl1
Z7sBaFn0jsMMG6LChpr0uNGZ5burvCuTmP/CiRh4OJyLX+2KZQcyJlPEONZ4r/k+hAx5Vgh9T+dG
YxupyRaB4V99d2/Wr7+RHofbG/vlJNDYk/a7PBOWHSk4ZKcnigolmNrtbhNEkmxV6+e3EXB6Eg34
c4dmDTTZVkF9KU0mhe5t/y3ZSF8mugOLxYxOEDQ9MiwEBqEBvXR39bvUr/DeX47I5pnJEV/Wy5PL
N1ui2gaClFSDTW9RLfp2RG3b9D9LnSQX150NUf62R+5lqMhZfnJBq3Clpp7aduB+oSLA2s7f0P0a
RRhwwAagw6Zal+xcVriLJYdCs9iNU267iZuiVXawTHZyE/6go7q8y6WN9uGUt/P5sGFqLsHQlJT0
WxQEZmh0AZp/bag1UsPm+JeKiETUSEVJeQme73YP5TVgmbvr9b8oIoimebmaabexvTfw5y4tIPWm
rLizLvvgZZXurEjhtZAjgN38A1h6kmTthtzkAr8Xl8KH5ZYPFcvl19s6WWw551HApgUw7PKf0huh
eK5MBLaGAsp3HSvMoKXgeak+YUD/h1V+ksY3wYUyJ8v+qvxMnV3mtNVkJk3j6gucDvym/0CXOO1N
jHq9i9mXgdVBHJ3baE82HD/eFwruJgsUuGaAl8K/7hyfb231fOgEzFZzc+133S14zgd44d6cAdMz
u4yhCMzXI5GwFQqOc5UkkJ7oUVUPC661J3hBQgVx19fEw4OGH8BdBnMXGcnGqaXC0X1QoXXe5+58
NSnVKTPVTN/gpxO+qkR3GwZlm9q+JxLTo2FBmbUqKAVywszadLBc6tvGA0y2t5hPQo7heS7Jf7AW
LzSRAZtxG6wn7gaY5WT49AL4SIUQDFuaBmlbWmpVYAQv5nlq3to1ExRssHnuz7tEnxZEbvz28GL0
rX0l93EqjGiGoUPZSUq3aGSPovL+2iR1WVPAdP5Ll89Poji0xIaXbbVBxvJlCNO+Y/NHvqYC+SVI
iimpeV+4dRoh2aWy+nifccqHOAykc+7iJyOMo0fVZiJZ5olnY+PzilNkQQdEo1B1tfbxmzn3mc68
oTHY7G96UgLZftadP1h7t2zQchg/ouv1ph/36OebRvi+6pyImfTX1VDmx1qKn+CZAwt9eAbjrQ+J
KhlSlhiDRVMUf7Sh/sV4ePAXzqE3kmwG5xDrx+8fuS3xS6cYX2p7geEcuywbxllwnnUj3xNc8liP
ah/1lqofaRZzXRkYuc79A6prnCTd+Mr0buv1dZGG/zVXq6igNe1D2s7r2UwayuuMZRdKghdvJtoR
VsjfsCZn4PdhG09cxDDbX/WmiBSwRLE+KtzmniEZRVWAghnaIp1njBizs/QRVJRVRt4Rn8iZVYS/
ePNZY4I0XDTBSgaAOTo+x6yXqt16FifJBtKTF4bKJJtFcYICmSoyfj8JxSz6O0w7Cks1NEwlAa+i
zZzMsCWFmKFIC7D33TrkZZGzGBmRcda76aQKrwt2P1xN4AWqUkcmNuB73g4KA526NQRUHOINV85K
xoyAU42apvGoglHWUR86pQhWK2zDe2c6bI08zdoWZmbCUcJy1s2VFs/SQAvn5rsMljK8jGmiD0qh
eCu5hAvIbyrpRp98FNykwJ3Gy+aAeKMhrMjErb9CXx9MyMizfWwGzDbVCvCqUBvddN7P5jARTTNC
aURNMX8Hu22a1d6YKg8lAqNIwgD8tfjhnk1FxHbupY38/Vr0YYN72L6BHUYt/Lvu34uhvAVBNZyE
rAfB+HJ2XYzvbW7615YO5C3ZAAKRIlN1xoQ70S3pd+eLqHCDj6e0F39N54h+3w2BSjcjVn42UNPx
8viyxT63nFusQI5fDnB1SpzPyuI3x+LkrGdDI9Hr7ERGT22ZuPo0R194fpXgtS9Is6C+rXZLtc+Y
ITRD4ymmct6seBRxH3N20kLINBMF6+7isPhAhaKNmFJ9aBRnrY/oO+zc2qNmd+/sKW7HgZV+f7kR
uuvdheZssSASO92p+5tfxOxTjoiWzoLsyCzznDsjgEI816uv7bcgUTsbwGypVt3fA1K56i/pMQaQ
4gwwweGUeNu7MWuw7gsXooSrpDCtsUiiSRxouyBqmh8mMYk8MSDT3tFcCiuk1+aibdIVr1ltTZ0O
gOoVk5zbh2T5YgWOHWo0+GmKSQ9jhGb14g3JgJO7ZXRsvODuGRuhhwDheQq+1H6Vz/5DnzkDCYCW
uGMkuVjeF/ymKS0UHlT82c5kC6Kje08pTPEgpJM3YQPBgs24dCf7qYTJOu4PmbM87ZIudBtBV0aN
5rcPDPCO1luMfsKjDkkUptPWWI1XSmVM8UlKocQsKBxTtVupmbFBgyhOZJtPXdvsa4SlcaWskF+t
2K7AwInfdnYKkBKRCa6MsTbyHRTQkwRWXPrSOjy4NtXDPzu7Dir7HnCaz6zouCQ68AIF8b2V898o
PbPiDyxcbQKHCls/KH5+6A71rM5Q0mXmRTnKnEg/QPGxXOzt5FD0fghF/87udcYIsDgnBIUrwwFy
CumpCqiLvgAhhHtFcYymILHsOwD3mbYRmnS8keA2V+E7a67yXDBIYzV663gOeh8zXCWnDye2bMiW
U1X5ctUiJqSfblsWdfWxCjLtz5WLZAHQYJgvnQ0zpJTigwW8Zhb5Pu0njw29cH0haNdPy1Ts9fEy
gKDmczXZuihz+D+OwJv7ap6ZxorQcOtA9NqXEohF/RITdUyDXpf9lofieh9jU66KM/Lvl1eiEX4A
mxK8Pxin7uD4ugpShQdJjGNZqm29KBW3OjRvdJrwtQV6QM2IEXqdOwOTjBaBih56cdGPznPQQoD2
GllVQaD9qyq4aB2P/ojbj1KOLey1YzdvTlt+9A4kjZZ7zSTmQS4Vvy0qVME3qX8tNGFm7HJik0WY
/zGJ4AXjetAQmsWJlUQtpnMkZNDRgFiDRVSEnJ6QJ0UOly8FGp9pOZCo3QfKv+4EsRlC16DiKugD
blARYnTi+dZe5vAaQq6D311aQ/gExvkzVqbYb1orGR2KCKbJ3D9C4vHWazgI9npOnjoIEYJgwveM
X22GL98ypQycOk2yeXMNwrZoHxz5tqZWyuiuC2UhZ89nU5Z4Metuski4nGmh/mxSpCyMTnPjaSCp
FX0TQY+etV7w7uNxWUK4lpIIOH3oNkwBAvLYBfuSA4/C1Gu4z+hMPuErTdtbP0okIHmRl74yQl9U
qO15+pIz3EA36HvKYEz81itYpCFV17NfXj7suQ8a+JukFhCZkTizv8dh4l/ULpovdVMW6/PvHZ/4
Nld+oULh8TLmo64jxltTpUBZBtSucQtOZ6Ikc/r+7MPmk8VDVOlqwY12QYy4FPjUojOYOgfgfPpQ
iT6dgmd899IqSZvW9czFroY9+YzSfkcMljqFfaWms2jNmjCsBPXn0LsFY82ngbTI9NWcOACSk84P
cRrRH/CuqVvDCWWDGURVYDxz9ocHX266P3ak9Vj+NbVC7eZFWEUBAKPItbFQ6KKypP7mpi+1yGqs
TcQfWejjTGh6XR6FS4p15UR8pQUGUu+U2JZGSIUgsQWDrpkUf23D8iJDwNtw8D7IOiNseuImI3aN
S/6PE4W46SwF8NdKyyFwzSwUI1SJy7j3/t7wr7AvR6nb0+5H1JxHoy7OY45SMHEP2P/zegvn/Nx9
imD1/sFPRUEQSfCEDv0fQNr8KQMkmyLQz7OOZ+TLkjghCPAsQSoAJkB7q+Y6ttnqJ/STs8vx7W7I
Nfy47GcBcJrlfxaMMWQf9VqhUQSPvnqEpwDe5e5odEB7neqq40mdBGvR/85Z6k6BmlO6Y9gcuAB8
cMLfHcpBrRE7Di2lJ45BCk3tIFOzthhLrlPzOPIiTGElLr5oxmBmxenqbsKepmnzUTfO7mqzjoF3
yaNLmlvkwjYU3t8XzCiOrrF1//ZkfNa/NBp+/7NCt8vzGc0WLutq+oV6CR2tYFCsWo4lxjEiMKFE
Q7Z2kKNaoBDuNNpHDzy8c3lCtF6tlemYvWMScu3MZtZc4My47K3PO1WwENRQ27itjqCBGwBW8mhX
lc8FVm6XumNFOHPXUxQ8k8utPdeaWzjsb6KWOkDHwQGYTmw1Nk2G1+Hb+Z0iZT9a1Vlw+SMj+3Ek
jkj6auhNlWR/tvsdYupzpwK3wtxpqQa4gVEWET2EjNL3dOUsxbIt/UQvaEy1+x25JD+wHCAUpI3/
rjgMxPSaP/pL6Q1oBMWfNe/WcJmE/6FiyaBpD3HqON1nFry03cwhS1C1tSUcep+DrpkwVXqfScUs
Nvvw2y3B68AomaZmcjqeJ+p6Fmo3V3UnBSNlVysbShKtoaDkrI6rYDBKqWoBvLGeJ3Pru1WJbSmv
SLGkBoT12JyTCDrLxW7gfEtlU8ZLF8Gt7lAg5Ar2f8/8+MYa0Myrvbo/4a5AyfQrSpWHx5ysTp4y
gtwWPQXZM5iBFKiw2of0vUdltIJOfVqotkmnJCerkH+mEb2n0yqFjwGYJ92eXHXDaV2bA17b7eWF
RaWJgYNuQrjGn9Pv0DrLl/0FokGE3KZrXNq7kxsABz8kUEPnt/kkN3gTBPnOv7+pU2sxpkkCyqf5
FdQOr7GsSS132ZIgAa6X68LXqK01OqZ5hxdVFbeojTCLrQbIT97sk3vtc5ERWP5MLQHXxRrfYPgF
YeiccJJLyrKaqeanuVz2Kh8pKmWvwkx+cyFbww5amLOJyQoLf2DiqvI5jE7xjVfO83v4JEfHhj9T
ttRZvKwQgFP1IvOsZGtjhwMYB/+cObj+TZWuOLiV0NUjuTF88/aHHg6J5LkQO1lsi/zCOaW6pWDl
WhJoh4PF4w04l8+c381JvcdB+EwX5PtvgoiBczZSwEmbPZFkk33TFGP9R+fbg81PCN06wgiZxhiE
AKpiHLmRWD5x9nQESud5kkP3LDSP2OtSTWWXE7H1By3zB75o3FfIv2rZBjuCJBpLE+oXvnJjRAWJ
vUaU69T3fKTMYYiHxI6/FnaQWXxKvwrkahsHt2UmM9ip9E3VkAruDHZJNciNZ5OLcCkmtUg81PrH
hooI1EwSneYF2N9jB+NR5dwSCQ1pKo5eRVw2vk57/Rh19uJVYfG/xNkpSc3tME9fe/SsyI7rNOCx
RcokEZe5Q2A1ZlBr+eksgTF+IxxoDG/B0Q+jJlHPaBBvvkjmjd8wKz2hl1etbR4YZjgVLbcVPy3E
0/nuSJnRQUwh0PwtfDo9RRe2jsJ2yOVjtf4B5WheY2E79+VpZsGm6n8weXI4Car6MIBqGPRdMvKL
B2EboaEfTEFM1ab8BaXInaDr7SLv43/hXBPgmtoEowhHpc10lZiYCkq3OwsZEn9e+zHuQDum1LpX
ou+VfEIx9/jRez6TURve1VhRzP/ojqloKTeh9kdSGixneojXxrBlweM5gBmMthR2gaU4r9RNHz1a
Fkz9At2XGxEfppwFhW/Xo4ep5FdkPynJdMNcFqlMY7fk2rblbpr8sywjggAGi7kW2ipYd9reAMir
fQTmvG5sNHZY61B9dbu1Fz8uwdK3h0kyTzMwvpFsty+X8ecCv1xrDWtysDnttUiux/flkXpBc8jU
S60H9YV11kabaFd3sSNMVOJlk5LP1fC+hJXhqj5Qe0hQn8VK62/D+Ut2AtVGcIbVezQZ5NpC6/AA
70z6HBj/jVIYXxP32PJco092Jft6KX6ajbcqao6Lk1sOFkYlUKLUIVxTSDxABkIXMQCOYJHUp0eg
lblku6jmoYmCqHDhOmwSQRW6Sh0VV34Ywd+fpvrSMJfeGhkoSnXoXf1HrjIs29ttGvW1cwBRwIzR
pRFMSqwPq0k32k/OW7b+eDaXDSLZDyRwzc5h0sUxjyoP+sO/dPhpWAaDYqelwjoAeSgowGBHTXI9
zdyXUBt8lvaHQUri3/N5JdZpRBJ8KyUWeqIRbT8YZIsNSXIFS8MNnmYfPFeCEb/C544JiBcqknxm
NpjV+NXfp1pT+JPnvxhV16wTu/0bZswJolJZlbRGKP6eSzwjN4GJSEYuPw04CECryHKKn7lbIvHB
+UldNgom1P70FDJK0jGOsr0jHKggsR20rBbX5SqDz8wzzVRB1/0DZTR8Qr3AsYvpkfE9XtuCbEQT
U75Dosj3bLgRg6kjFRjC//FuzAOGykcFZhhiqepcc8bie//Hx5EsDz/9YgGrKVNvJQeeYvw/lEDQ
ccB1do3IP3b4ItbOSmL8Wouot3MgHXUpIIDZc05DYI35bYnBqPqmLqQ1Wb1CqPkkfMjDIY7/Zqqe
Jh4eAhS3t9UBlsa867n0sY+0AXRrzpUJsMAhzhrjhWhfgvaH0Y7sDSN5RaSmy+Igu+y5v1ZzycBz
rCWQjZLQeBOGrlvmvfPM5TyWMDYMznK7gga6l7p5zkkPuQTnyzUDn8pv3HkhPp3EgcwmL75T9Y6c
DnpDwoVJKodQRG8PJS2cdz0npq9KR96wVlpDvcTqRCGzkg+0Z5Zf/CJ8FDoWoY4p4fhV6VB492ka
0/DAna6u4Pz9KC4UG8zZ+p7aRMiUB13NasFpX5Ilsep8he63f7p6q1C/NVaa29aDDpv39w5mpRwB
4rcnX2TwRcHQNveJI/XVcTAJKcTbitjyOINnsWP9yl8T5Pcs11w6p3u/mLedVpYgBnCPBhAv+5wv
OnN2htpPUmqpqvLvM6i0tYxzEK0YRfcSxFgC5GqrG+/f0U1ph59FGUfcs5A32y/YjPkzhphd0adw
rSyKRlDOKu+U7O0TttfmvpE01IVb6wrsw6L25pbL1AB4Sq0wjqxOb8ndAnG8xOkeb6OLKCWaWUe9
TS1AtNgLAPkwRLqolUz2xRVYqSSKzbXCJCvtiZVYlMx0ZLcrAY6oghQNLsTqSWG/AWjLWMZkeaeW
FMKA6i57czNB7qqHtFU/NvJfq49zVdJ1Ky3kcOgxwyVdKxx1J0AByn3fLFOpsK7FXqkH03e6hXvK
N7Ld+0T9c0SGuivvGab5BMRfhiRVfYdDKTfo2uP5ovmHksdQdN5ZJyM/yNfshk/bsaXOZ/cGcXVz
bUMoICcYY5387CeBLCZ3We93Zx06GT2FGmMXMyyYrRyJBDYK6uHjkH/6jgQZY6hW+7uLYpYx9Crb
MEdaX8oDSbSHNgAW0yKVaPIGyW/Sva03MyQp8XRGbW8Aivyzh8w6ezxdMGxDcNlDUzgU6ZYkPma7
vduyCiPIK4Cv0izNkKoh+uMgD4nVn5SG2gWm8vjYMYrctbmIEczxud4UCQ2mvrx8P5KeKjaPmnEY
w5UC+IBzxAv9b5g2qIm8bOn3h4M02UGlGJGqbwwGSkE3EppBMhUisdDrZme7f4osf+cpbuVErNFN
IMoP5Ig+tC84XOvm8QH3RdFjUuvjzmzFjh8iVAkV3nWF+81l1vnXAqunjb1p/RyoEo+NYWpIYTp9
8Ucdc51XGO6GA0cC9AciRubG4KvLHQdVZlQgWzCwDUCHKNZxLE+onLIXEvvWaDefdg9N+baKoHjl
JhNRmG+3dqwHpnFX75wtxqCEy6FQeiCmvCAK/cAvgeOILQ6ufkl31kbNuo7eOXD5K0xmeVownRQ2
+xg/RyvwwCXmv/s6AJdq8DBh3a6wGBFdceJZh7LV/JlWOxvFQ7fAfP/QEjtbj9Y1cHGoVlr3EnHm
yrK/OllpIyISBnun15P6J/S9OZFLu5ZTIFIYNU8Dqu3DUbe2o0qwbc/TO9W3mfNo9BpKXEOVPp6k
/XpMCEJpbK7//rH+/Q6LJyL//9WaCAbcIqa/m36Y9sHAP0cpsTY/U8eP/m/MH8y4YAzE8dPjoOZD
dtctTatKfyWVmNNe+qO5JRzGQGvP1HyUXzPT85sKDP1uLsElVPO07ZGqkdJRU9STNt1sTF2WYdcl
jVWhu3aH2Fk8iTBp5szac9XwBWIND95WIRNs3AzqIGGXOARSxtaH89ZsNmZ4II1owMcfO4KUZADN
Dd9OOsYiU4wl+X5ZQsJCTPf86qweNNRbhM/pWZ1USBk488u9gTvpm+RiQ6Ky9e5HvcGiDsnTkz/g
2mNE+49M8CchZoFHARfAIZkfpTN4milR6koQPw3u59FhWS7zWJ/ZkZ13NMpgPlr9QQJNiWXXCG5t
KOXtBIrDdUBYo39r+WUDnZ+7xUeM2GCv2rA0u+j01Dcb6nRxkQLt56zBh4fgJyvUnAclq92mT8C1
/Jn4Q3iHEG0YmsIYMYPqRICxOp/V1RkhIjkPeCYSDYIsmItvWMNbzP/6hWosyeDqfIiNa+mPlU3F
H1kG1UhlBYnhrfpnfJT3VbCN5YVsd+x6Hmp54zM61q1z9eMWO+EBOqpXnQ4eJUKlyBI2kZWtrsQb
tPnI17Pbg48BMuQJ6kU5gEm5aJE2C9HMH0cTydBsgDHZS6Kdcy9s3GEfQn4tt7XT/0Nphx0gj6IM
fw5t5goNEzIB/tsMCkyjGdZ2Wd5vl3PxjsBh6r24voODj5erieiwh1gjxwKzMzJszp2jdUj1TusS
+e/xEbtjEMr4S3OM8aUhzpaOchO10CBHpJEGoesXJGRlx9/DD6KtWPVSSODvJWMtfA9Yxf0MVdfc
rR+m26HbXuuaS6VsOGGUovLziWBpitPc8SHEvpO++jrryTMrb1CdU0LY0LSMyfsKtwd6PRGhNZDd
CeQU2gvcbIut8Jatecr76mPWaFbQ5VyjMITJmSjHEbP6IQfXBRFuiX2uEhLqJ/BBgaD50MZbI1lr
/TZczSz5tnYVJPHHraK1YR8EhG2C41jXgZpzayChIc7Vam0BshdBNXovTttmYBbb5ZaFgQIZQMzt
US5a6RAit1S10yzC1X59p2wyBgCv/k8x57nlh8unlHRU1G7Iq0kHh5e8sjoKGYQsQdm8NgLXmaVB
vNRxlLUOO/pSsI7EErFAJ32mAtPhvThkpCThTtPaSm65hBGNrk8i0RhQlo7ilF2OWR7B2Qn0wTCq
uIZm2RqvSu68fH/TWZBFuZFik4R7a49cTUxnEd0KWh6o9H0obxtTvOpjBsp0QH0oAccGAhVDNYzJ
/3e3O7V1kjQaURVUaQqAAFaqIoVtWRmRhrIrLFiQNi21BhDjbXsPfq3cgwLXBwEtnBqD5+jghKur
Y07EzEm5XmUq9AYnqA43bBkk2eaCbUpn/iccoq+DG6Spha9UrTIPI/ifOxh5VIv1pMspKFVoCzXy
vIArwiEK8BxkP/k3HM3GubifVuTuFIjy/vZWqi+ZA/eajbBf7HF5sCUq1t8OSomqXNKU54vN02AA
9jb/59ckJCIJztPvsQQ2/1Makn52scu0BsvdEBiv2uljBCWpHlGrVLHRZGWMUvsDpG2msMrMIwme
6XemXw/xsjXO1o5NYqttMkb2RZ4u0k3Cf7HeGcKanr/W1AaWYBeiZrnrVsT8zM1P1WXW4wtvg2Fk
Tdv5FBi5vxjOXVJmiKEuEi+XqlEUhB7hUy/88auYmBCXfceExALyyktTXTZXpUxXLHo59/TKskSA
S96KlJnVZ2E8DkC45/7WNZJAOgKnPiqw5VPX5jatiyf9q72YEIbqWYvNe+ZWRVERspyChuvx7Zwz
qePFDHi+BKqLXOYpX2iKQit8z5sBZn98VU/OPpd+fi1KOKupRUbLSCzVc12oFQwU7pgv7sDHa3Aj
W7MTNIBgguW41catBgWXHrKR/4zTDC3X+uoqsSGocpzHaU0CiJ3yGTEWVgXPYRdlaz4KyvtE+V5f
MU7KW1QxP+qpbJlq/IT6eLnITBcepuwJRvOD+nqlB4kS1zM+XjoXqqL019G6ddt87Z463Z2gDydv
jWRIDtRXBql8zjw0KC5YmGU93wC1PKPEr9OJI8NyhkyZuDbHcjBVTB8w0RMZrtxsEVn6/GbIeg01
vpivLpmMU2l3i14mCQWQHgYjTYqTElbDZgg9y/HAQiCU2QLPgofX+nI71W5S01+R0GC22AEqXrtO
znxYUfyfEC3rSEPbbQvbgXSfrsG1x8u/D5sZnH8v98J6+g7AdO3YBmD7PM/grXeIWh/bz7F0svlP
9K+8W5XXbKWx8qpRt5YPjyFr+cNB9zjiYNZOsUe4j3phxeZqnw82lBfFkx8MkB+yxK58NJwLP8rX
zf6bOu9cJhzakrbOKuJ1rqB86z2dTDff+JPrjprFjmqFt4izy3E93pFgo5w7IgdIpRVdso3EWTR0
KLNCWCUgju0y63t1gCxeDZwgHqY0jQoKbcK0gCp7W9qS7a/yhXN5SQFchbi3qbROlxVCLSIL75Jt
Rwzk4WDUO6njGKCZBFfbKkOWDdterBN5lUphgru3KBEQsSdK43LExjBpPN0aOuKP/G5LtshexoxI
wrK6zQfTPy5ht31rXfETPlih0ycZs6TpQPoksztioCdU73m3bkWbtOOpr2hxsgQA5KchTyK7VSky
QE7FAH9qgpQFJfMmi8ZiHZpzlHldwdhwPbTPHNRUC/xldA/3XprWgm50YxFC82UvlCoAS33Ljugs
0JbGW561wsPtIzdssnZSkgYd4K1PW4vzzOe9kHFCzgtyK5hr3vkQKW/JQZiSCz0vLoOUqefqQ07X
C6ky+lDqvWCUs8mf93ZWSFGfH6yF8vEe7Oq3iajWJkYgBRf2xEnYoMJB/QzZWh1gKlq+h/Hz3A3g
gMWOg2fZtTogIY0hEEtZQk9uLaH+5o4AAIVRJagbW6GqJEXXdDOgVqtsi1wbJ1LQGeMguotC6MwM
O3Wm9+YYQAMPcj4ke1WCAHKLNp91nSjNcp/2wugoixAmZ5B2eQcIXKQXoaTjCcyzDNlJ1Aq6p/8A
KTpv4gVInJ2sxGG9IiDoBFISjxNXwpog+vTk/1kQSiRpMtRQMCBFfdQFGvGaD20/3imfR7v/Fesq
LJVvpPudefnTHddUjpYRuCY+KrkrbhiQaPcV1wG3yurp3wb6bYtzmtBaEFAcXo6RVDejuEpyhvAB
cKLigDsE6GjOwRj1l5yb9CanRXe1GbthZ5Vh4Vt2VsCSKYXMm8fow5NWjAYihFJlfy/dxjuRdSmT
7OAF7qcilOZCfzmmjps3KKruEwllyOno5YODBJ/Sv1hCO1pVHlrgMB0ozj87TJ+ptgNmXfsx1rtB
1kXOZdAp+WSnexpTxRkUAiec3zy9fQ46ApM1xlY/Vk7iiDD2nRT2hqAksapN4OVO1FXyCWjFh6PX
rSXuzWO1gF6eZi80NMqluEJqlPA4gszxoMjOMiyDjkLbaSYif68QWVAnf2D2z5PHu2VaugxcKA6V
klm158A85jCQTbG8sFxM8IdFJzAGw+tFaHxW3poFX4uEYGhfTOT1jkGe0Mz70tldSQ/3Mfmdq1Bn
St7lAc9fiKxiB8vcmVAAKNCADN9ewez1TjhRUnFj/Ytcua34MvJM6SZbDolw+9oM0kxpOiltSLVZ
3ZebNugBVoKdcdkLHYKkJaTBFo9U21f24qBhlMj2NzMGKJNJ3uGmmBGiF+Qd/JMSSrho5fd3ShHr
mrpmeRr4uNlaV0VTk35nPHe4eVT4LZtzarSStVbrcC0aNDHBpgCCDdoDcQaOd619tRLCLSkIr2kd
NXrmywMaNsaYC55EITSYgUF0NthlGcyWb00b3CftujclFbrvXPZIQpNSwb6U2oBtP7V/blDIfBYt
EWI66zCh/DSa2Kfc5P389+nbP5RyL9GCpo4XDEs91fIEahGTh2l1gShIMQWq9C2J5+5P3fbu4t1R
R97LyEY8xW0/iX5UZnmjDCEPvDjhbLn8S6ZxVBwW4A/zIwOXVR0niyQD5LgwBKhYda+cFr4b03Y2
rmGwpzl2dmPeX75I2i65TQIYwoCKJiZO4PEZV+p0Qt5OrM0UGraeIXHgFxBgeABpLGPI+PJO8Idz
lsMfPGiR5d+u97XFeBySeUbzQSW2vKrF5ETAYyXHGhu3Q3mCppEWgtZadTHP4hkSmRLVduxz57ps
Bxg2Gr4pF8nf3iorttoOk5loV5ir8eq/uOKWf4rYF4s7E+bofZ4VgXe0+tIR8t+u2ed51bUYo2jC
EaPn96pR9YOkQuw2Q8qU/kULVpjTw5ErWfjjxZAbj0RMDpGAYSbeqmrlDnU33pRhJQMwqKht3gRQ
dLvI/a0s95NXskZc7ZGAm5TGE+xMNLpi3ngvrwYSXXSYg7gJaiwWJlABctdWyS9yolVNQusVSsvR
t4G6amvfp0Lv8U6+JDXjakm6s54SC8mfwOQn7XBjFNh8dk9KacqNhPxOexemZI8jjX8/j8ovfhvE
XCxUxDiuXljwN8hIIpYlw8Ka+it8K4vySaUW3ju/GhOAxZKMbJtbTArTIX4hIrhI9/XRjCYEg9vN
L1Ng2ANqblcA7ngGSXA8pw20nFVuPV8DjBtte13+gF1hWIaBJNcZGYzQiY2l8LkBaLpFhpaVdsFT
MR7XqJlyIFvCZvWamR9uZdfiAVicthW3MAtPSG5NFp0OpwFUuNT3Wi0KiXmXMlHNJJIdiRFiaFgj
2SmnNcwZHxSfQ6bZipSVMK907zpvlU+C52EXSZoSYWxnCAC2PifaJiaNKXNB+gnpbn7U8KLtKrmL
kZCAmwe7QKjUrAmKPaArYc6mdYuwINYmS6cDPX3LUnw9gGFm2n45Pupegpdx+G+hY2acsMWZwMRw
8Gm+96jTZSVVVeCK8dhKtBIcv9O2ze9jLxdrHl3meDeHEt+vajtDLxj7vqr16tvTeWKAQR3+uEJW
LqwVuzj9Shc8p7/f0Ix2SDMf2X0QVUXOltA0Dnd5U8yeoYP4xY6t7NBvgj92iedSgv5hhy6Xr8VJ
LHMFU61hr4mAFGZ2eTeUs0ZkuuMXoVQarxtE2atoHSjSyNExd4wih85rOEV+IAV/kCa+TkW+uVlE
j7tc7WU8L1eLaL030BLgVg52iZYfKuYbDXYSmUas3kdSU3QiHA7tJcYOdg44XZOGKH7VTDp9tVud
iIdTePJr7t1UiHSl/m5jw20TjFryVqor4tPLO+wQdTz6Xij6fKGW4YVI9R+5bLyjzwHgMll7H3YK
1yqePRjgxTZM/w68UrUq0tbqUlgpKe45Er/Y+l4NDKucBViaagCCscWmZ+KLm6OqqsdeecWREVYD
skRRxUaKVFRa9h0DO1AjkA0o2mQoIorVvUTywcPf1tD4NY+4QEDdg8wG2ikHNEOMX4AkGkswraSC
nBf811hRxgxRVwXXS3m3dYETKYKfQe2y9hS8qTzRZLjjQmmiKxx4EnuQz8QrwnjvegAlV62ZefWG
TkBUQt5Mb/Wr5EvkjB6A1ItyzMnr4fVj0xNUUpvK47o8obiyPMg+igZx9wM5XZD1xQTiQLiHm4FJ
4Vgo4lTYOk2A9dzRAbh42bAWDXdiaJMiDW4Htg42mg81yhzdq3OZL32rMpQwANDfHKP/l0p9tSe2
kG7K53KO6e8cUuoco6YIxq4onqPY5o55KpumXKyDgQ94K0LkxI1arBUkfOVAxEJEDLRLh15+pBZY
OfvQVuEqg0BrDxiDdXUdhMjpilnvBGSlOLLpnTz7pC5N0n0ReyUBI9OBDse5H0XLgNBEJZOo7Ua4
EnOWygyN3YbpSHi9C5hdemdJQ9jR8YpznVCSpCNKX+ouOdOWYDhhBOJvRWBecF1tr/ypb1HJBegC
xQTVzpiWsJ+zrhf9TQSuVFka4xCIZc9U4HRlku3pOAyMjFyvZxqnUute92NGEeB8wgjTsrGLfIrY
x0cJq23Am/QT9wY6KSiPXboxXVBU3o20AVpbH7b4ym4nFj2VlKyPAcpZq+rjYjzkNNYGCjkTbc0S
hagk16lnuzI9FYdiE00K3WmJbUI4Jr9U5KInvJy65wV2pjEVcDfIKJ6jOc3W8OdVzli7IpzxDI52
8i+Zx+MnI/wmV1ksFwBkLi2Jem1mN2hD7C/0rldEl1ODZ70BOJxJ19t4ZwkCcsfCwl7uoPqZJrL3
ph1rFyF7VFuoI+tZNwycA9xim6+hAn8NG2Z8dhMnx6FL7pK68u75jRp/KGB4P0RzvWI1WE/6pq05
vYRa8c2vAM4ZyVP+nqiKXuMQyCbntB/rTpXnxf1dQvMwMudjFPDnpKtrd2N7n91HOqrAOvRGqnjm
Mwn+nfTdRL4K99IUaqouiaBIjCkZ1gvmA3yPe/9HHUu9h8NQ+NXnhM948PvgCkyYukIChwONaj9S
ha4F3rR3NFvp05rRYL8lFpm2+5YZ0lRarDVNR9NKOKgDGFNHtYzFRbtaRhVeNZ72XsEKHcw++bMj
lZz7/P3wj/E76FRt1fcHyPESW7mrR4aT+QZq8VeRkXyE5h3Y1L6qt1JhLRExAgcaaRRpjIXXVobZ
CaLaHHdypTwGl5Ju/azrpLpWBPjXi4881yL56+mNN9Ci5MjNIwUq7m7wVagW148Jm75ZJH27tClo
JqndJ7GPSlpB8JRqTe5C+rIQpGeS9icwm8ZF8cTft9wjHsUu8Z46x7yCIVTKbZYXzZ+TNHq9kKkX
eFDPmepKALr4XjoT0mxVTdWWlu0v5g81GvarS3GVH1wMO+GJ4E2BnRxUzccmPCZIngUQVQN17Epn
JqMkKfOJ95lz0V8TG4dysOXhXIo9Y9M4srmr/jAHqCV3o0KTseMGrvHc21nWyoqmdvItM3ad1SVq
J8ubxtJdMeg7dNCWq5XQ3cywJxIj/Sfe5QhdcyPTSldNxu3Y9m0yKVvbDWdPN1ubNvlPck/Jwwd9
0QlGRYdblxMQoFY00LeqtLmMEFtqbCpEQ/GfbaHRP2nLiwr3370RZg1OR8xqlh6uEI14X2go6Hn5
Q6vFt/tbYqabw1oivfnsMxgdLMv3dLZ7sazEM4eNCYjZjWmPxl9NIo+j4GFEJui1KJNsKBdYCmxS
WTNFL7avbUdE+Osjk4zgahmDu0E8AdT1s3mCLE63A1QDZW25ys5/ykYk/akpsXC2mOtasrYPg5Yr
RtYxhF2OgYV6vKPaEoQd+Hg18hdmHlKCQ0auVTGAY9zon6ZH7lPxgbARJvQPVf0/UBXqBozVCEGL
7eeUDjGebCXhSROMORTNrPZD0M65pJeV6gCpaIcJPi+oVktqOAz674Msaqq+jZikLs5tRvxOkCvV
fjD9MtNGVbpSzdEoz9o3X77Y7CY3dluqQ+CaMp7mhETPq/2JZltzgF1ARzJAGZ6n4q4q3gpfK9L2
AKtMZacPVrDdZczKEOgv5RO7KzRJODWSqK+1TKa2ZZBx5nFlzbdRetmHZIj7egVu+c5iCGHoqcBc
Hd9eEtiLbSs5EeNYvjumHTocYK9S3O/l1QAmrOQiU2N2CMPLNvfoFWxOZRj7aXTJYNLd4Lqmzibf
GRdJYyhdYvCA2+BG/1z87mXOyLpRzfKf3Vyk8ZKyeiUKqg+UhQjZ3w13CTm8p2spsngGCv6a8+b/
+CWtzqprc+cmTAKm4dDx7pba6ugPL+kS9wq8Cf9pFMpVoSeyG/hwYlANaokzblJhob80y4cv/bz2
ReryfFTpNF3VPBD0mgci+r9crz1zQ/MU5WT4bNm9q8RZeWz4ImaXj/9eHXICZKTK932aweBFRGdm
+LRgFgUNAGbd3TMjpHI1vIt1XmJP6MVqqEkvpw2fNDGp3TWOyp+4mwIB8xFLrNt9ouz5QGAjLop6
ZnOXXQLtQlPIcAAbEKpGhPx0DXjpJS5UGZjFFe8QOIASHY0G7oMuqkWXPNazidg7tVPZEzdd0mdr
iklPw4vKsMc5aSwaLY8BMCHQN8xqqsTcXE8cweRreeSIctm3VveA5c80OavjiW61zcA4NL9+ogyE
f7ULuIkQpYSJnfk6HXq2VlnMXm+Z85n428RmxY9DkY5I4xfiPzjDHgeR1qr8TS52EKsERxEyIx3M
JHpGbDJNYTGW+PYImoklSDoKpUyQWOmrjniQoYYhgFLxo/npMROIMI8Qma8+8yvEEftfpulLbKSg
7srNxzqPcHVctAyWYee7VeQjNuffx/vroqrQVCZgbEben7vM8E7msrh/3DF59Th7kzR+6uH/gFx4
sHycPCaPZxB5CQDb1R5z8daTBZnI69W4xQscFP+7l9Ftcc9SE7I/lrDt94dLZBOTASS8bc+tU6IQ
n1aqjnUEiMjrNsUNcCXKNgPU3QiOy0qmQLdOhErnqgHI4624hUkFXXGTnbvrcKGN/3eE1fc+0qfB
NnQBn3Mhu/WGOnyHHpaV4owg23Owo4jSaEXVRgxrm8wgTjPZqqxdlcJvF2Dm3YyP32LdHftSIEY4
FREiQ6kaC+W3gGocrwAO3VE5URTpLzvntigHGRa/i5hCpSqDKTDGytDChQIvuduE/yVb/Cwy7I8g
rPLIMtHFjJ0yqlc2QGKl/LRi1TTrzkCK2l2v+5TRWditW6JdLYFhSYphlbRr870qVbv6R4yPfXpK
yj0PeyOBmnBG3QqZvKOBS2QN8q5lCukdnDfXMWPHQ8RSJ0NWCEB2Sf+v/DLPsoXrGRYbRwEs9ZUb
NgzoT6W3O2NLdO+rxMqkv6VFpweu0KDJqJY+rZiJT7jR1IMwhNe/WKmxuqWAPEgHmb0N6jRwt2Ts
NEK2F9j8LYzmHsqFdDa+scFwPQ9ll0TvzTci2EoWubEcahTWwASbHDj37/eN6PDVkqncYPSfPo6x
IzPk5wKOIenz5SopIb99hrF1MbLuHljBdbSsU6AbR6iSVGMOzL127yM9A5JZP5Tpd+brEPqXAIcE
iMjbukxYVBqpm6OuJm3QY59Eso7l0yy2yeSLsrlAviUgkj7ipFrVBPHJLLb+jkZjuAvURZGIw5QD
p67O5hbH5Tvaxj8b/oVU9t2N070nYQJ/0TfRacGUC7Bo7IDKW/GAAOGfHLknFsWIsxOlUTzdUgqN
d5+NozfpnHGAyyWUUBv7x5XcmOr/0uOw8RJ1ecWcmqK8xctzbW+FMaH6meZYxuxqdqgQGnhGTyuc
MDSJEwOd0FxgNmaLo4/UsD5tPZo9ebdt7sC7wBD6lButA+HSUXL1ygS/tkPkoCZVvce6TGM1hmaC
znIMdaLExcYXZlCZYweCY0esDxB0enQC/CDjYtk32qH1PhXJmtXFS3Ycr2Vm8eAN7Q9utUhchVTA
hQE0dYwMix8QK5xNXYGRbGRZ+CWiT0wEa3dB1L0NCHZ36XGFw60LK1T0eGr0AGRGEADyb+AU0Wes
g8salnM0M3GaXRIOjU053UO7wpT0MWyRmrO4qV2BsxU8jU5Dsk5wv43NC/YuCuL9PPaxsza8Wyh9
WFDaP+e7CvHzfr3Pb/BqVa8Fjfx3FybRLBqqp/0jZgfYVKSPDu/5yAfZ2bw5dAUv2XHc4M9LuRgm
fuvyeUXRUUlsKnomB4Ghb0cHrbeZ5Ux+i3Z0YfKYV62WtsDXG9aXoHrUVjL7wmH2kAEfAu7OippF
BN4/iQqy/g1Wuhz1JxJbvbswJmWNPqTcIEAN5dPUEPOllMjTCbt1S2RUdw027+uEHzy97om2Tb0U
heEnoz4cDlLPPdarOEMO8+E/Fq8IO6m3wnzGbb6+9zljrJ9WOVWKg7yHq9/ajzJEvxrbo/ZKVxUJ
Dh8bGpAC7uXBq6aoEQw5AovoreBVEbD4oY0hmM22Ap1MDLYmWiw5MIjda/xZ0oQp3+25kNkkf/jX
oR0hG0xhEM47tRHtvQvh5RL3GTD62bDf/HYq+1e0GAFcH2+4r9H0guTIHaVckmWUzJvQJu2fTPEu
ei28WIVzNYTaLJVcUIDBJIftjhVfbEQkag+wR5/8ZBhwS+uN1Uon483dl4mvgM9YJiQ0OWGT1Bqm
DZxJMHP0BF/Kg2uaaydjvYa27HpTUADDEHeTzy5F2AArxJaqeiYPLezcBqNFTGWtWC4GhTceFj3Z
28KoYm/61QXE+WZDs6+YqLKKj5EIBEbTd+khdgGezzGKYqgU2UxzEbFzu1C+G0dJaGhTABmB9N5e
+mWrGD420w8fQB6H2fYq93cVoLRJz9Ub2vQbIg8nMgjYQwRw1tbvRQvssChdsmRyXHSLb9nTrOwV
mLwZPQAozNvhoo2uSH4etie4FN5ycuq8vv/U58xI0NRUXsS/fsg+hHHRCbuZQCZkUCn0prL0LXHL
RG1wm/pyVibLYxQtAHsN+auXsUulttFUIIJhFSl04cJ9c5u4ZO1GxwVP8YxD3fd4dxQLDY1GRfIu
/VXHVFuVmgR269mue/yeeg1VJTebaUnZk6lKhmFEc8sjhZ7Zk5t12pe9A+UOfq+DjTV1Z8TN2f7T
vw+gRIqm0R29m+gO9k2H+90f/cxXNqYwx8eBowycLvUM2OZdECzWDIRyKgd058T0HFNlim+E9/39
00/Q9Srf7ZeMnDlpZhWvze9rwa9WqudXXylv21fQ+NEBDVYJr5sRl5HkKNTjI7prmK0YqTszy4QD
ZyDsHLaoCHhDjPEy9QYTE6UZmWADqeoy0G70YnGd7Y+sG6DSezhAr+Y+n6rozpdiDutMbgph6Gr1
6DScWWbyN3U3jNs2egW08JpR92fxvi3VVfSshih/XWMlab1v2/HJlf96DDHaAWvbyd7KjKk6Dzgg
mKvigxUFVtyB6psuyLwCRikeh0rlFVYG/zZ40QXqBPr/fqqbl49t/7pLaBjKd/RWOG2tXf8sAiqS
dGLpoVMGuxqjzUEA5HPVXwMbkhpS7no/wcatMOb5A1VPQSbfCXniuD+Oo6J3cjvk3N0NQzS1zvu8
s8zPa6IG3TjNDTmYNiGWjRXcIVy/yFMF/Ty3pQ6e77X6CIN4QK8adeox/BUq2vcHw4IAIpEP252q
X8pxjEGxTEGCD4Xz5bNlx5fmqviy6RePuBAoyP0pi9UznP2IeA9Sdha8GPMMZtE6xF/CFdXhs3Bn
3DD0CQ/+PxkApSV7kmw581V4xeUPA2aJ7UCHnEb7faoi5ix8UCAxHr2LiObroCiryMA1SaElOxUV
IwWeh1dult8ablIRPyxGPatDT/VeI+O5twZ/qvTZZnd4aEAPFI/1St49OeVUvDqRfRT8Uc2hrOCj
RqdTL33h0MRy744LDGOUhYs5i78qB0RFZJZlmjSuOpkDbDJrNiz9O6Y+Pn6aubO0FI7mhpDxnmm4
Oy+Z8L9LDJ3pAqXwPdmKtPXiyEoigFIxQvvepwcjgWllgbl/+JBtSVKGsE87EnLkOfjB8QTqSFS7
OUVUM6FPWDgzFSx1aO2DBimLwudEb00mQvNPuw7C9NIfJFzy4mRg36fU8jPEGREZ6uelYy5CT3r+
1MKXQenl8PUetwZTE5sHhkhn0Pr8BGBbw3GJbFDKFS2iknP5d1bWsC1ssWDwaFctVhVnJkQ5yXzM
oRYEEAyDYdR4W7y44IWHx9OPkvnAm+KLpi9yFNFZ7W40mRWSlwDB0BPpp6u2TwEK1QlZUe//KWpJ
npPW3ewy9jCEktZARwvqvNDfdaTnHTt8F2bmKHGX85IS8JqTlx4Gz81IAg/1JcNN0OioZoLmdvBC
eUVERW92RjkjDYL0lrPFyuVLn46sDHqPXrzTWaaPV7pfK/s/HDScsD+3zJr2S143VFEI9j/SoA9h
lMJKtNEgj4WECg8tUzgZMNuWAUpnIYACinsTpIqU13//1QTNcFPUEPr9ZPHAkDEjoCG9vNd3po+w
/Oz9WqN3JkRWaUOKBHq+zgwD6ckNN1YsK9ZJS2BSJ/v/sPfPBWFAjJJcNC3UJlff1XnIqwjXdaLO
yLW+yEW6uIk+IikSY1fRpkDCBGoTho+KejkYVPtDrnlbW4HHJ9OlN7HJkeEH7U7M78mfmQBUml/K
hZfaZWY8NlpPpR2q5PAv6uLPI2zl3LtrPQuod6/7iWPSvBDf5utKaOfd7mq6C5TXCm7L3+RpwGj7
mKs5KoIC+8m5ev9V30X0ebnnH2h4rM7rsSVX1ivG6wpMDK6FazdBplIrFdv0KoWiV2xqm4MPfaAp
wh25/jq7Fj/hKl/4nolvNg6j2hGozlLKdVISG72pTE/8jZjtaDv+dZEUF4rKOV4ba9KyaHms3pic
+jIDMpId+MpzoF4n+lMtzRpEg+0hn2lowlK1Hu3FPJAp8xIMhNBwnlHYsSbsIT/j5Fo/9MIYyDB4
xoRu37VLqxsFH3TvLkw0ilVYGqy2o8eeQNlEvkbOmkpwnIIrGi9NbpvB3UYydzLGhPE916KLLecE
dOFxBnURQY4BTdmhxbWh6eJLFveix1eA2fU8JwzAcAM+pIgIyd5hM6SOCQnJGpnUs2uIX8B38HeD
4ilnln0MinBgRPz+VTEXU4SqSr0eerL92Tg3UU+9pBAsgIVnjOT4zzKr59Vm+LupW7GJ6ed6EAaT
MAqvwhhuP5nfwBtJthhNjNDM2HHbyEILGG9osmebTWXGn8tgtMnH8aH6LRzLFUYJaePCDiaJX/V7
PTgVo3TCG1wjisO9rgDa1K0Dth8XtUznaAsGkrXUXyvJZ/a52jcLAvM9iRpt8XY7+yF7GGaRj40M
7YHaXNA2wL447GY9TKqY8xQ/lNTtcY7aCPrhwQaNZ8kaL0CSp1ykRKDEtxF7ozHYdIcsAz3/M+Z5
10bQVuwmm6UVzKhJFRHKabDpq+wuUKK13utTOesgUOpJvmM+zPKZai/7f1WgbgCqN/+G936cCHQ6
7dX3kYK2gm9tHzfvB0YHEc7LHbtZKP0VCz9LMUg7RCQ1mnPOvN57JgEk8IZVSOOFDWmId9pIA6/j
HvIgNgVpIzwpoowifeunH3g4nZGAvUziTiPMSzPVmuN/D5auhKUt6jWFGiEQGqZBnGItHFnM6iBe
2/Ocdr1zcPpN2q1JkHOTlClzCAn/3zVzShpQKcvfNa+yLO6QHcRiuFA8fxz6QNo3TnXpPmQ5J7ZT
RIzKbcscemL5LrYzmQYs0KK5kAE60EJqyj+tmY7/qz5Mh4q9PEfIZNV6UkZrTZOybi1mQqGfzZJG
0Nv5icZ9gw//CbjV/k5OcfRuoFdwRt87A8QQUQY/s+uopMYTBHjZDBoadeeAg5CBFjSaEkLr0MI7
f6/cNrCXoon5Q3mjF1vawQTaocGH8Kq38Tq3m6v/BvHcPhOHmJhtf+uKEmgv8dRRuKARYN9E9nM3
u2PDZPdBIcFIQL48AOcacEZXnMVbJ2ema6n8GtlQOcxrk9R9CAnN3aPQWNlFPH3xhA0mBXPYSKrr
0ei29rZrf0IF7LC++eUMRirsTwiS0mNS/4fLiLwFxTbS+is///a65eUqbZQVxbZacJMpjnA4c5N0
9tYhGxnmEdo0+DCD8qIL/9Td0NZ/1ArVtEp9bxtmCEICk+gJo36KfCFwE7NCZGETJE/NGxUu1+Lf
inP51jXXZ9b98UtgfJyEJZRn1F5ifRv2wiZBpKG5UP8aZ9eWAUUBHHJCeL+gRXWSxerLCzLDjAJM
ScSqvGtJel5yIqycUpNRfDijPi5GTojKmN2MNP6cOuZ4boKA6HGjt8/T13ZLaOafU86Sa3+0ct8K
+Zcr4wCbFp9Gaf37OYpRE/bGdTYB8MMu5xAJwMPN7mSF9bcB9y7tg9NADkn+RdEGca0DpNpwicMs
KLF1pN5otMtAFyRceKNDcKzDLAhTCPt8+5gEcqx6m+g1bPg0u4JqOjq+Ek20J8hBNxJ8Nolqy3m7
Ky1nVNcwOyq+BYwERwbl9I1Uk5CJlkeXMv2dncshhGk6+6VPZq60pDYs6w8IzRQIqUdBDGcS9zZL
Ocm4bCC4/KHrlsscbyGz7zWXCbTbaPkUpYHBZnTjxlkNeQnzaXicIzgm8Rh7B/tvrh/JnclbMAO5
r1xiBJ88j3LR9AAa1hyloPTqhJ03NNPKL1PuRRVSZ5KsWDeO1cBA2hR6qOQ9it+NXVuFeTIvX/xA
Jeev/RbZNiJGcdeRTZKvPNTzsUpoqOyJRR5fBCIGwhkZtBObTdVl2JfRMqxz9OWNZ/4BIE/SUilN
7JX8ss9XXr5UdI8hzgxJSAwVy3EBCxyXZkOkMMu8W06ZiLpf6Asqn8qqzN+YMTDGpy+ydKO0L3Eu
rpUd5tOA1WDO7HTR5SIPH2QChnuirxZMroH+QzR3HGvZg2BZHZss2hVfx5OxNAiDmdpVuiNRCXsJ
n6hGCpolzKxzzFrWlLb5CYEYT1RczsD8PyyAra28TJz2T/SN1kJbvoOScwdHgPI3/Obnmmim9JVb
miWIwjvB05CFHeqZj2WbNpo3IgI6wi5/8q3AkUm+KjFyemSaeGnW8QX0nNAfdQKDYycgk1cKBH7N
fl+1BMcxcWgO0qKftaUGCF18vNHq8sYUKZ1uFr1dFmIP9leH66BfoKfyGYl/4GrFyppjv3U1NZLX
BEyjLPqy1mB7z/0BMoT3saUf0fgi5MvUPVbRhxubMY1o5t9V3h09vn9ewMc9edGpxvLRA00fCGq/
bznIeHRGa/z/1bqtDJN+2g88uAwQGsec07/cLdzxyNQiklHKcuXidbsikEQkiyvupaO03Y623V1r
A9b6yA8PkUGS759izkviio/7biE2g1S3VP3JzSeky9B/p1RsVsuaXmkZdeMuj2nh3nb26U5mVS6c
k9iLfik6oa0fyb4mOx9VbKR6lSevqyoPnVUYdnOo34AhRy3X9Ndp/3+tjM5kVQ7EYaaN/spjmAP5
YDiVautA0/blWHjgIQdpT7PIp12nhRH2ZvZEiiC+ttpR/REkk4SIkUNENLGBMJjcqD5vZH8/QK4j
m3bhUeH92I1L4zxAjyQ1lJY5zyAUK/mdA/gMAstNT2jKoGnhcPRJiaLuZmQf1K5VQVD+o72+ajyu
iF23Ye9zxpFNUC7B1Hgl5OeTYPFLwnM9JLAWgo0eHqt8NYzEMddD8zaomteVo7CsJo/dkOizDFi5
Puh4rczqWu86E+Oldx7mz0wd7UClFUvURuaItzlm95mHroyKYy/klnqa6TpZHuodFaK0tAyMo9K+
vkJlbGApw1V+VYBKtfxAVkTW0K6jjyJuY6gO/95w2dyKBnUnZaoSHK3m5dLJNbnGtpnC1wdBDPIL
w0fs/MrFIXSIq/VpscvKta0BhCGRvtSHUJiM9PYUhPofj0WLLGVs2s3AqBStxe7hbhpk+YcxHyJc
etcSVlc9y64/DJo4etIx+wNpOww/SY1DgA/yksM2Ru5Y5axiQk9xVZhC+Gd5sJhCKR+fIBZfEX+0
nwIqDAm6nz4Sbp1Rny4u87mvB7sioqaKMpG7xqYpWfsaIVn56G+5lzL/UDobmI3qZXnQQn8OmtSV
W2MQl9K7imDlrGhtM9U7Ygt58oIZCqctPxJKys+MPQfi8TlUxuS2/pXvYaPL1DckYnfitFvb+H3k
962UtvffWcmG023eVKe4oXi1u1WTbLsoQSn3vEo3JpnpCdTrUkvet8OBE44DpQTbRVu6VCXqIYDE
bnegGdKiXqRKOsdHI3XlHKmKHmEj8un2f6Oa/SMmfdfgZoZgSltoYcVj7PRpPNg2q5FTfNr/lbfI
CjRsM9AX/FPwn35J4qo9M9AjrFccPkc8vQQKHWCtZpo8lvR3rdawb05bFbC8F/JdVpp3vwI9iKmt
0rH9ad9exK2473+fWhx8AxR8zAF62VhJYWc5LGrslgkGW31rFj+q1W5RJKYD3djaZJc53GzvuVCU
PlZN4HiM+Fpl+/kGETwYzlDzqUdlHN7JkwOT9r4c0hmmugDAgASry29QPw8V6bSoTnkP/JY8s9BP
MbK5INnPEVaSAPeb6BRHnhVfEiXS7NbknvIdHKKMKX6jRQSKBQoMMnD3bh1gxXKvYoZddZHzGyiE
fj9NtP3RQOc7+rxo7I/MSkJbeRcdp5E8f/ugPipO/FxEC26a6gMxZJ4N/QPxbdKueOjVpRirU3J/
PINpQxMf4B7lhqkCt54pdM3Ob0wnXTrWoTa6jXFJnxROMqZv+LKBcINU6oxaiK/Os276+WgIzkzV
nHUCMzquKCEIS562tUFpdkJNNAleXR0v0FfIEN/m+9gHcePU9xN+YzeF9lfQgaGJkCqC4EZKct9R
6mrvvtyOBCXrEj6JqG+pqqgFXQ5X33JJCU7ToKIIKScpRhiLkeIANfMNXpNHvfYMjubze/oNABOz
Wm7KK4kRKY5tzFmoztd3iS94vZJF8yC1gZh0155rVnr08er1F79mbNtXz7uZtZwqbg7oYwNGA/AN
WEiaYW22u+ZabV5oUMCC/rXAN4XlXHRVhFbv/3zGMZgOsXsojMaPZmtvsLhaBLd9Rs5gMLle7IWP
7WLzTA/jgAyH92J/dG1xtZlezwUCArek8PmhcQvx4V5GVcK/xmWx19L8ust0OD75Dvj39q+u2RIN
QozST+TJE8fXffUTnCJDNxRcNGrHHA0fZQGLljDsP550Vj623YK/4k8V+7A432Ks3SBtn5slMlj4
On1TIR0oFEygLjwM1TyNYNdjYLLdKm4IEuQTfOvcL/t+58tloQwHi35IcXI0/nymBdf8kswV73ud
t0HZnYTQU0VyqicU6Mc2h1GhygkLrIPYWG7aNmqTb+33yhYr6OSUqMAhXYkPW8dx5+Z22y0KeMQk
ssNMsM7ezi9kGd9QTHvRWtEKBYkzV8KJTaInAc2RA28vVzFim6ed3GC1yajn1f13GhGlfUe4g0yR
1Cu8PmVsD4wPnHJ+ymtl2bj4Lu5PrPQKRyl1eJMVOwnC9QNcVkuU28wiEYiAbPjHmNO9KrA14iym
ChkyfE2sHdZ7WNlt+P1VFs+RcE6CXgv5zsCCzdKTMdo2HjcihLlKBUoNJeFJMvkXqtUqWYMWuW56
4XoI1tXvRFqSuo0QcyVUccbZE50uW7O//yN9QpSKnhYl/7VfXUWZ6O8MdAxl1/yVg1uOsKPZPish
6Gya1PC+Fz4qucA5pcPi7IkhweeL4EILp4OZ5TTO+FAwxfb+ZbJg+USnO/b6LWuZTehkYeGXMa3C
GXEH7BrWdrywXOayOa5TRJdGDclcrRS3pcr2bs+292DNj7tfev/UI4UCrPG0Q3WmVPX3jld8hGsU
YlOV9wvpEdlHOPMZh/I3PO6MLipkuHTmb/mV2Xe6OKjXrzgs5uvZX8/uP0FMZGQEWsDMJ0pGhX/t
er9ba4UE94NKQoxbcMS13EovLrx6j1eIY3ST9M9nHMASV3NsbDdBlJ0Mcdx6y3WuLzzAn6mLxXmP
/rKdRatRmdsmX1349Oo8lJZpNM9y0Y/9x2LTJVOOBYi/YaeHlpBX0PIYEc5pKo/pgPambazeMwx5
UpDauim6fDQSiZv1lcWECHgy/QPzjmnxBiHvo6brJwKYCs7jtmbl72pkHPdDxoJ4MNxsyExAoUix
JoJzYPMumqwj8sKiR9D1igdUEReBhvVzS66SmCM9ozocvdgZBFxBrpmYJOUHiYt4G6CeK44okcBz
6ehL1GBNa8TLJ33zDKfK+oReDhH1fc6jEC3kmNtvP9jcGeRagZlvJeM7lqBzEPbB6QMal2nkLLng
NMpzCcttN4IVDXV0Ap215WBobTNdxram4NaCX/CNIZ6FWFXAN1ckzWRpHfqAJwY6O0DIVUlWzLay
rXyzJXLBs/8ssL1iZh3bz85dB+9LE+H0iGky/m1VL5n1CsrY1/wnINT7UhTDnBbo9EyAK3wjbF4A
Ps9+qCY95vvHKTROJynsA1Fs15m+oQVjPHLgITC6S54IUohJWa/loULswe/8Rq9nS6YWJna9stre
/g0cIWGWJLc7fI105a+nFZEmySiEPye3AUDsfnZo2xwCmKSP+7fygXgZ5qxC55cQw21WZwcUTq8b
cjT9RL4XNNo+N6QWXJaG8JJd6KRa3VEDlzg7B/HxbqLuV3PZ4P7OI4sUm9DHq1yxPjNKL2s+3K4N
bvg5aDcv8OVa7uSBk8zpaYbVUZOEgsXMHJyTkBJso+ocGCwxhKXmdJYjiLd3VP7onsNFlnJtepgb
O7e4EVQe8LSwKr/+aPg5HHsRHWR+E9aSkVteGkB4Cshx8lhP/GKJ459YYiQMrDDgvVSqA7aUnQrT
NHkmFlD8qYIuLk0wouq+UaAVuj3r5nz0wYweOGRj3Q+oEG1kRL2/7yZPvzYoFEkRX0CJy1+XwAmu
A4XKwYfVw0LA9Z6yW+w8HOFRRCypND3wWv5JraaWnzWVveLoM9w8CghhUoMM8NN90q5UTPyJGu77
DZOgQcZI5Zrzdt7OPffhy2N43HSX62GbVkaZ1DwcIsHs+C6wMT5MWfSDQqQmkzuJ0yjvRn+wXb3x
DOPcf7Y2PrBjBLoxKv+DTEwZ8wv9BtxtXKxcSp7U94A/YPy034GVXQREO1q3WS/k+RgVBvPWJAqs
Q00oByPidLicdJnooq63gMfUA1s2yYRxYnoatGdW12WV6+Y5skvI6Hk1x2QllA0ItD0RCi/1RnjY
BBrTiNqdfn3CD90TZkjagstjs+DfgWvRyK2+rvw8/xZyt/7VJmrlqRHsEYte+VriajSV6OCb77+H
HPdroQysP4l+RMsUbidRtlsT18XiBQaN5kXU3+IWarp14I6MDkIignUJpSi8paHUE2NDUIcHmlzN
Eprc5778Yjw6SmNqOZRSVOOaSxPVkHXj1R5Guk/93gsS6TmFBQmE0/qLWb20XqZ5dkgCSteDcwoQ
pm0GQrhgfLYfH6uVBPKngdTmEHqyENV/AdtvYtpxnw9GBNCnvWxXgwLnn22bT/dTM3VgJyHwHosH
hJo/TZJILZvYIXrq5wdNCnBPTVtBHyWMNzVWIDhhb2Rhq6b+n8mZDtyzfhQZsKDITF1qhiP6LcUd
ioArSYLsUgoGGtZkwwoBzB/Ql4mwmxSRTMUyZ/AWau1z51iT7UgjiwqoKrd8bs+DcUFOeNd0LXF4
KDvYjwtx5Y7gGObWa8RidI3nMKu6cho8YkfxXqXGXV8GX/hOXA2Ahwi0Ov51H1+12wJubA2VuMKX
506hMnRS6P00Z81Urjzy2PEZEUxe8S1yXct0w6udtpt2bAm0er22tY6d65mxa53Ko2vF9+prirrN
GLrA0T2Ckdy8G4tLU0jTqVQCkiNhbjSCGrCnuvW+cU0IUEWbMmTNMt7DDs8DOHMObgY/tVxvcBip
EXwB2f4RGD9kAwLT/GnHlzGB8r2ju6XtfvU4lC7ob7V18jU141xVQY2eFLKoBX6EHAI6mrMswV4V
zvprJqXWXZSpwGyroDxAbnqaveLF1dIN0iqVTKPo3dWvXes85HbRY8b1KqwGtuymIw3xtgNlShRR
2Pmgi8Gxjsn1mjjHqaW134WO6XG1W+hsmbFLzwxqDpXZvB4iQp//vagMr7vzI2ng2Yv1bLRrgUy2
OqIWkId09jJAvNqBhe/PbSZHlD8XkcMHyrlbo+Ma2jmHmxX78rgRwZufSnee+t4G3IM+kO4MBYEx
Ye7LorGb6Tj/VoGNFb+Cz/SSAPx1paEHXu0Xlz+VwsIOPLbj+0Vsaenv3QkuvCxMpdIaKBbJwBFc
TfNhNPnZ/ZvskOXKT2he9YiwuFIIelLIeyq73kFkqokO4ySE1QYcfrE+kaqvG9W5JqYWH9uDRlbX
rQpJCMoDf1TwtyCkYAggYzzEBBhaZKbzhJnBatCbXfLlgLbjdaSzlbilDmyBU8mRa1La1XkUukps
rWtOXxEDv/4tU/q3WrahZzUhas6n22gqvnY5H6HXRt1iq8vkSiTNzP+rLF8P5Dv2dpLsPIluq7Ss
QMI+Alg3RqlnuZDlyRQwXzN6UxhegOyAOiF/tLc2WYZWHfztwJjs98HJRLw4WUs/ROZDWxIlp6pE
mKMrbd+YKimVup7dekU0OyltK6qCt0Kt8tbbgFKGcoEVu0HqXAIu+eyU4+m3xHcJZM7iTNP3bBGU
vX3f4BIVfJV1dRa4S07FTTEqrZTz1LRFrn0/mIGnSZGRxFIzOXWWvrTh8eT4eqAxOJZi5dG8IDP1
hkZhbtCD8wjTiBD+Yf5zjiVJq2sUuETstE5NsHeUihP12Q3B/eQHtbmiKAXHm+gPpulZqxew8zWT
kuLvMd0bUAfctZ/XcnJl6qa+ZIMTuZS8EtsWcTYQBg1YVOcKXBSIoNz0E2tZB/AZ/w09PxDJJXgq
m2Q3BU+zy3r3xe+Z2Dw7OkSJ93mEVLLgrTXlr/n4tZvxeN4Yv6j6XW8cX/9FNqa9bohUFj9tvDj7
VKbYbw0d4h1vrP8OmI7ILh/DHsd+5mHTmPhjO3XVFLHBLgFhIKghpmYLVEYG/xWuO8B6tC6oI2mp
CMtDQl3cDGRCVxEXAERWafB2FOIPJEeVJ5Wonk1xaHNElWIk2kRyJHU/HAX8u16H1tNo9T2gk7wC
eVfl8UfBHqsiO+DfxiO7tHs5yGgYVwaG7dwvIA1qN5JlIC6gefyq1QF4JIMBsNnDk6VG8dYMq8ji
kX7fZI/HiY7tfF2x0ftdB7uTcsTJqMcFCT2D+HNnv+bjZNJhuuVdFmFOHyZDKr/dEaRuzHJodnIR
+shRKXw4iF+rUzsKT68BbbEFolEByKiQ903U7e3luVsNHqch/KGlYs4zhkavB66OblF44TQY+vt2
UAb7K+XQ4RH2038pakC/ta//pfRTwVrMnUumBCCigAaHmxkez3BXfrX9v6hr6jwBFVlI92V+Gi+t
Acc2x6umtT55Do7JhZmulo86F8TOVpMcQDUFI4Rk1k3m4U2a91ZuuYh/jCIoGp1JNMOPonBzeJOF
+xEnKXO28bDZgHRLS/DNqnkOTqr46TcMRdV8pBm4fV6mkpBZhH7+5yppDx0bdaSo/Ax1sHuhKjpR
fNZgzIWIkc9g5UlCgavK8szCkjf1uUMDvXmGfNDV008vdZK3cSgP2+A8IHVCVfNQlEwYfCVgRzrP
OHyjCl6ArYA3mRtKAr16KoyWdTTdgJ28AyKlxPNug9wrW22H1GCpdb2RElr4jafxgRauLqjCRWdp
GgeLfveSKLEikGGUeIzOVAzX37YJCO3dF1nGYvlFu5Z4r7yaD9FuyiufkZhk7lZduEc2D1LYC8e4
M72HprOzUGhwnMYfPytp96UvcyUXOESL0JQtWhzSP1jgyyECo04vjvi5NCh1kroC8difhMsAzEEx
8uQWPzumeFQ1jyBvH5V6NpwTw6smv/ChZzcnclaOgwH10k/39JvklxZN8EEpu2Vn8K7g3EHtJfn/
XNSxXEDW1iai++7xXR6FwonYei5uaez9Meuf2yaCUEvOfuce9/kG2gHx0lKC+qwCDYQ0LqKeRRZ2
btr1SD2ROj4ILvY42JygzM8XicDnaH1TURnRp+eCy9nFbofQWFUH/hrvqvVZCkkJs+P7ziWMFTDI
MY0qSto/dgZk0fKl9PYl1u2dcr3/i7oHb8rswbZWYFUp78CVCNFFtq7pqTvUVpZ5wEyGqxWk7wCo
wsJaqSgCFQRn7zOW53hZe4BbTHoQEosfZrkEexuE+kU9zNGxB66ORmmE7MQBWc9QdAszatC3yPbY
aMNktYhpXytyu5erZu5g1rYPw9oJ8Zbdk4S7oRmbFM+EiWWSZtsc4SzIrxDk6Q5bqXCmeDdpGQuP
OpbwOcBm9aTtetJXPE6lGfdzatd0ovQYw6or6BI4+yUoCsEIcj5ZNJ9+o8QUc8xCTwgeJcU97pCJ
IEkR57neHxxxX0SV6V7113nRl+LyUqmGaZkqfUQHPzgokZp0zaKxtIvx8KgPfJPLu9eYQQyFNWGe
sygHSoIKbCP6bJPm09f6gXiXcvEiDMRPSZ80WnhNxFxginiojFLgRXNU2NxxIU3uEGrM30RfVOMu
GVulu9Z8+ZR2Oi0ZX+wxp3F+2eIrA8XVhrB08IqMQSjwcY7l+M9QCrZ93Jw7vAujwKFyzGfpSUY6
dfqu0NxUN8vryagKZ30R6I7xWrsk/ag+vSTNlY6ge3oVUMtLX9gJ5tXuCU7m6LWfkgRlSHqQFqqv
gWDm5lzxkE1BcobkwVtw1XD2E1dOTMcOYWpGkHy3nKJntpwEeCPi+b1wdcMVxQ4j2u/qNBgXMLs6
OfjtrYH81j5ijW6AduF9IYIa3yEqSQjlbPPFWSfG7P/ML7O4YVGpEjcidJABdm+Bjf3q1sZShaFT
MW3Zy61+RMM/LOIoadlZ0wGVG93+VPpv20BweJqaTPp7hxR/T4LSdhl8bl6G92aMxZnEYhVlcJRN
KbX4myETfW+IwPJ7v7ZrJi2f57Y2T69NRpulQ2EJhNVdmO/LTSe0AxnraZNIULWw9vl6IOE12/vX
6vsmFw4uBecBzqK2r0XOTJjFeniNRgzGZXEpPmLQPM4LE00jxPx0HvUzhZjvLqZIGXe6km4gUSQE
h2VILbmhjoVGATO5hqZqfQduR8kC80bnmMwgA3JSHuxotEJJiOnvPtSSn/TK2vWQIc9kpOyO6fuh
1vwGobQT5lSxofrNN655rNXtM1IKj5sRHNVwF6asK2Fk9gvo4NOnTq64hpXYQvwUea0/zfVnj1T3
+pNycHx+KZk6JINu/T2rmycpZvRnqNVc+e0Ygeu4QdlS4ssXA5V/kcQmryJaLTnB4I/RjrRXMr+u
k4MtN5PswAvyfv53KVRSG+jSPPQRLOlVZ1uy0yDpJwj6vjWQs8AgJfx8QsIrdOsHldO+NySZwUqU
GCzTIX8FgGGL6ko7ZEHt7OUe40EW8kSWbrX329nLMhWs3OgpCNZTBWn2MIPT75NOa+txEws8lZEj
5gyDkZB4525rKPXmIyMZ6DRHAtO0M87ktvk8D0iQoF+xfP/4XqRiKXmy6983Zifq3Vuon/LUQNhF
qTM7RxlXcMCedr4Qgyoz2mpDAC8oYDVEGnDnEc7yXdZ6xoggX2ZTZYolL5fOw2t62R2NkDI2qDo2
SIvDHnhFLIwBaE7AIkLJNjiI1I1ndtseEQCrGIs4XHl72DLaj6163i8y9KMAwjm38baRmzPogqIB
tNRh6CJ+vRWMSu3BxCPx4H618pbjXau1T6lYRcuB34aLrLYuyR5rfMpMQwLPEIm19mGO5Egq/h44
1WgND9ZPzZz8QCPP90/ZrgocfY9pNJIZ1sC4HKQcj9I7g4nI6RB+FKO01V8hvDYRVM2U5FXCZ0Mb
ELQJ+nhp0jwCZJwgfu1i1W45zAcwsZ2/Q6ioB9eyIpG4roWgsEqzBfXQUczf688DD3pX4BqYjvNw
At8AuKKw32hrtHG1c9r4AUgIzHzHU9RQSb1dM27+ej/BEJglH5CeXJD13v7mnJK/1R0gnRKUsINu
YqQv0Gm6HT/4TV1aapXj0IDyvvsay3OZ0vEu4yLFQF0OJrpjPWMIoFEAyDf/K0QQU3CYqzfNbzy9
DaXMWM4LPtZkLANeTPefNN3p9CBpxol4DQABrnPdpu83isQrI+ZeO/ZfiGLdgjy8fjpJ5jkBgXsS
4L0hjTybonTD165qJQbnhgnFXn349ugG2LNeQr/NyfdfBUtpaq/T9JlShWiQ2Ci+VEx8PDqJaijC
y6WUcqhlp20JWYPpjJ+ZrCghaT9nbaxoQfrQAOlj9QVspc/k+tD2wTON8UEuA7D4hyvcSv37q3SF
5H9Awa5d67QGsPjNLFP474j3y5ruG6udeqYSUMuq08Z0aq9nam9WihEcIFQ8Pg84sQN0IaFkCfJ+
klD+y8pGINVypgdyO2AtOBNWYIOctQ1num/Jm6I17JZYJgYIobzsGhI1I/xnvjprD1E5PVU8io0c
mZXR9USQ22PDzOlyjbXAa0FyhA8n/WlA8I3ZRt4gLDHjTn1Yt1E4t6DB1+dm8ohYYOrSQNxgMxTY
a+c4jOXeC2u7sJtX3Q1Szm8WqbR9bgCb2jt1oYpXDlzb5Och2CohOL9u84r4andapykTafSVCB38
VEfN73em/JvO0TdQfeDHvb4PvKC6fbPZG6h9Ayzfu0/cbbrsZBwslWIPcO+/NeNYajIr15MLD3lO
f2dCHuW+9iF2/1iGDC9jup3ZgVxiDqOTyT+h+nq2i8HKKOpvXFbWul10p7sfHxAoyEfo7jhdwBtC
tegE+Dktwjy6BgIeUHnZixiNKJY8pIbaYr1U9jC29lCzBNf6ui9BqxFQe8FR4Z/BKpPKk2KcKQ4H
TCFxaUxWzPq6WL4yQX19CvQsIpB5FnD4EzEiII6vy/A+52IQK6v3q/qpNyDRQYAvIyLm5AFTSL3N
zYrTNSqcmwUwKaZf0Pa6JNoTSDh0O1N0JNeF1hKMXSPtln4jKqD+nw4iYO7jAs3MWQEFM7Z52aMh
Iyyrt7P2iORB84ZuepuJFCiRF9A24Hx+O/k6lnnSGXw0SYKVQw9oZeur80Vj55Cihoaryns1iytu
Xk1Zz+KJY0SoGONn3a/qjLpmnsAg/Rivt30gwRMPhmg3Afn8ZF5Bqy48WFtMHF5ewx8Gs5jnKTCi
MHG+TfyhlKfdQQTtrJV+vDN3MVyu+Fvm3TG5yJTvribJV1svvVGXbcivanCLWsG+hO5ztQjjY43V
jAM54J0OG1Q9vab/iczSRLj3QEk9k6O6xBMLh+4iMawx1wKpatZRoiUymYqaopwUBJqhNgu2ICch
hW2VXRGma9pGNn7c3KQO9h0ekvCCsfpvdnKVCOOFgYb1ncCRBgpLxOXmEOgO56YNVR2d1eNEY4Fg
Sx3mnQdOGT3JkhIBHr/AsS7HXh7TESCwY2tiP6RxkkJk8Q1H0ojdX8tEXM41Pkvl96Q1sj1fdL0h
S5135XIJO0dLBTQ8wamFzdhqy9FTpHqQQYGSvZmJE0vb6SIZY9k4zTKYa5sE2F1WvqaqpszK4d9w
ZhIcSGc+YC+R0y2aVjXjRvpUbspnxg/ICbTFGWMJKIhBlKv8juH9iRGIEQbrVR6KGuFbroAKIbVg
U8XQXXOg++7mZ/FW9DdD++ug+ByqzsmXyfz7ZFIX6v59/Bpo11x4btdLJILaJRyykINVlPjH5o+/
hOGm+As7ElZtuGSWfnRJ9Fe/D365iSyGdvjeQ9Dd2l7AHdup6J+kRFa2FysOp3N/RL5jgv04CXv9
xtQTI4k4etbI4VT9EJHCFopZfUJHeSVT6Dzw696fjvbVyfygp5Q4QSMEyScCDV1v6PrlZwnkS29g
9TLbE6A+/Tdd+IpSFyX61bEqxjoGgd7xII5cmgzktDhQ0U6eCo4fyCo5ZXlF5n7tn3PKUlbfUn9/
BXxZHlyB/vEmsdvHV4tiD8J7aNamLNSs9EgJcuUZ2pI2mAvDE4EObn1WBcM69AFLqePT3p/hMAuP
qHv0iNruVSnGJzc3nR9+MzWGseAR0IfCIgIeEUzcmdfl7EZnL5vwU0Bb1CjTJzBRkhTC/JpS/az2
GeAerYLBYRFpLWPw34Ox3XoA8o+175nnT4HZOoQzl39HH+7RXzPj+Q/aLfpQnzblqrE4VyjKXmx4
C5vg1dY+6EitHi59iJmXtCE3iEWohqqJ5XEsJoymqvEKviYJ7yxAike0BD5EEI4bnebZEByK6XLi
IVzN/AjQ2KAS125WgCbm05sQmvt57Wmh5hLMFpiGlMOUkjn1p6Jg8p3h1htLEDwsWxVH9hZXan4e
udhmbS3jJJMsKoFT0kKLEOpLr8bZdTJ2kpQF9n2ju2WTnA6lY8wWVE8QV3AD9gmkqzHgt2Qdixt8
8Kgt/Y/zJja+hx0QpM6HkdpiZXVCNGcV1mKRvHuMaodZ+Kmaa4JHU3i1DKI0rAiKdHW9Ix/Yxu0n
BD7XBobB9Zrgs8MXpyCBSMOb3eZCwvji6fSthXdiFtAHTKyYArCtZUHsA1NbciA9uGcTRX6iEzGy
ep0hkyx/bjvsEe7KximSmo2T+JS9+VH2O6JXG2/SWanmC+M2Zqt8y3RdYFZ/2J99JDpvIwhLWzRI
KK+ROQpIQNce2yPsy3C5LJfAdH+X8Y19SaLffNEdqMvk8jn3Zkf/v5sQipGzwwe9rOIjiGGlhrFH
541pWiqsic52OhCN+ho3iat8NrOVmw2E5IU9OUTTE02ClhT2HOv3QpUqsjz3uK+RAt5Of4UXW14q
9qphpc5yNrwaPtO7enix/3DzBuJIDGW0Fh2tMSFP4+mNycO2ZxurxWoaXC08Tsj14EW+9r4+XNJP
psjlrAPezD/PtShYhUE1SwiTNkHqHgqU6P2v4OGeovEdUXmSyQapMeIeHn8xRMELwINuOdoWYPxg
nVCGb2iN6ZRrGkchB6/2w5O3Y9AWK4SbUeqwLG3IbxzPoVl4LTUCUy9RtBfmlreRNfvlX9nHd6Si
cqvwMWFyo9FyJuvQDn9vSFeu0SGiyLZFkl5iooC+QnlH9PGyyqoJRhEPFWMQgs1NIjdRaEac6j/z
bsJvoHBiyRiZxkVi5ggVA+ke5UCBuu+UI4IoA1b7FGYO1x3fxd5uUp9s9CeGAoQixzXbpQD9jLql
ee2tEXyvNJh3cHEsi2gyc32eGv2WDho2wj+5fmz5yUBHj/wbDDx676YugFP9CjKduV8SMjr/voax
jWaDcDKLEsUg/zk4wJLQUVP56DK6KBTVYVle6vKC6pyaH6RP/I4eco6gtKFfLVLgLWKNiMwrnto/
IuCs5JLIqPMZKWJfT5PU3LbmU+uxTzU7zXBtB9O2YpXBpUTZOEq7X6mFdegoPJ60rb4v98Mcqr02
vpmzfyF/Dj+bgFBP+nqvgWNGyRVxMTDkSqEuTI5/QA9/TlPOzygJWsksq+O75JjzpuBCerqY3rYj
/vh2SF+YgVChqQjZdYUynkJEC4AQpGgfal05v2Cz50UbV3OJ2fjohoAMM8+9/ggUtDpBTkVNwp6w
ulf2MaU/wn76cczj4Veiy7Xh5C4XgJt1tyrClWo1N5IUqxqJPAgDVPKZUJRWSeE11LLj+Toip16D
7fnJNuq+jIC/3k6TlSLpI62JQ4XcT3ZiS9nqA9QQcre+06n8XIile58URx+IobIeeEp6rqKXtIo8
BHo+7VEy4oDxyJVMAUo54mhdFy45TNbuB+jXrF/sMOaIXTj5YsPMhjpx9hbQXVsK9/Wbz8RG94ld
05DggoPqsesLrXMRztfE0Hl6olcYs4c0vTW8fg2MbVf3dQ5RaEo0EXkAte/vzeCIeEr7JgHEEWO/
2Jsy/UqxceUi+jUqRcUNHSrJjuym7weI/VhZ2A4l1Aihgr2/9TcGyetZLLvaR4L/Tu47G/pCm4FB
EV+pwlTa1Wz5s4z7SG619VWuSMBtCVQ6BDCkbpkSv9RUOX995Dm3YKQZiZRD54twr+UNIUObrpB4
hGFGjLx9QD0CbgNHGQtmsa4kGyn5bhqpD+nVD6cTmjAz4R+AiiNeIoEFp7RXikWqsbhZSJ2dk5Bg
dFffKeKcng3/TseFGMZgGL9RQErTm/IQunZi5svANZJQal96uvcE2txgirHic8CKrqkubSfrriMS
Gov9EriU6nNqrOfO9NqzOMQuKx7WLn9Mq21cVXzuYa9XI8ICq75XVBOXLwqUUoGtlMCJAdj+4XyY
bA9yF+Znse9i0mh1MqgyJHL8lnzl26Sby8aXaeZxaASJia/YXnFIKhauwUqBeGpFs8gUuJgw1riE
AfIp+lrOkNscQbaFzsOLn/LurLKT+MY+TPqp3STb+vmsieqKPJJSSZpv2uIOMwDdx8mvTPal0D4N
VXbH8HSS1q1IrI/13HYHrJs3RLqV1dolpaAsfavVtVAtkQF2Nt3+nvMUrIYP5ugvkMXEn2OH6Uws
zUadxyT87H0CxtTErnQPqu6RqpepaC+Ao6S31t5mYs9W85vQL0WUhKEKs4V1NJNLaNy4RYwZJBbs
F00k37PgQl2WEos2USDD69dZurPAFOb/aVlg1f8YanW7MoipFMpqd6ZC3Xe7igWEFmVqda3nXPsc
7vfUQ7ZZdILHlZkR2NJZk5Zu8IWmFGTn1WWbQWoKKcMLYKuxSI3SvWVyhBjlLFHKXBx7a3PT6nAm
kRivkJKW82+PKe77ahufdIGtWk5zWmM45es6lMh79BO3ojbYLDXrcImKTjOrFJTpC+WIEUYyBbi2
awwWE1D2M4U/MDdVu4N1Cq/ohqvCdQwJ+xJ4BzKbOlrQww8eGmf1KKdEnu8PwNozIPsNYFSDOZUj
9/2pqJZeK2dUfb5G98qwBrIn98A2ypayLwI8DjXtZqdQY/Lddj47R3bS69prvji1onfKO4Z5NmEt
1tCqEfW0FDl13Q34fneXlu1wxaGOJz60XPfoYiZdct3tD3MMMoFFUKqGxdJZz8UG/2kID/dYZCvt
tJWyG+odaL/4RO1vg6XoSGuzxPr6N89ap7uNw2orgNut0d+hx4Ek0+pUko1qCPqZzoRgkiIl8ad8
9mEFkGrx3HZqAuYxH+Yuh4RfCSPAxeqNec3dH0mU7DwV8XRqlkQXhFUGl1EQKjMWT9DAN2qE5YUI
DRgF3EGte1AWrfzUj2x9LtVF7lQtUHR/GBWN3GGQKYFfCZmkKkUAd0HD77goNgn72OzWDzqU+uOr
MuYimevVPYsw1JMCBvLhwXV4+q8ZHTronmLqNzRY3KaiowFBnnj/o52a20H/Usx3O4BPYOmRagM9
LrUdTY96fLfFKCmdQQoIPKoSYmLDUk5oH2KG4ZBZpGdSqhYexh28JGp7VC8d+TLdMXxMG8JUcK3H
l7d4bF98si6l1KAhBv7qFPnGOQLAtF+kJfzlmaR4rsZAj0+21nVeosiGqnzM9w03lZHKIc4Vco9s
aDV/X7E++6SOfw9SwvnllgPxnPrhGcSqjEyw/8OsAgNYIGdm/4t9FIoNiy1LA5ZjTnn7cwqaMbLK
luB2aYaQ18vMQZNolkLsCBbArFkdbl5OCcJobpPGBBkB3uOQJqzgR13CNyzHvjcFX1RcIalyt0Br
5zff7PuqWr2Bno8Q3PP3jg00dxWVusv/mNDyyeEZxq6JpppHinkkNy1XuDnVti5f2hn3GOKtIvcI
Hld57KlHRsqs74q/ROjW3kb/Y7niDDZa7Aadm4ueuJN9wCrD3Jv4ykAdNwBop2EdYV8U1H/cc5uL
nf03A+g0awcMsFPEd+NGqS6MRJxZe3sC1yIe/azQy85WkzZF9mzun1AiXdMPH1dP9l3eHMnHoIdn
1CJedMtpe1ej1Zgl8DAjkdnUqgrkxRp2/Hxe63+B21Cjns2zsGk+BL8PKGYLT8zdI1xi/IT9bX/2
yElYxtcQsTPOeH36Iyxqgr0HQZZVd1yqws3OACJkw52KuIPQxK2X7D1Dcsqxo6BaDzHVrnrwYyxX
LLVChjzemha2FsZs+qJf6P1iiNpHB9IPdoyCtnEsRbXkjMNi8ZAj3TOGlmcNYcqblUc6hV7rPPwB
DKkR1CYiFSVlOvR2TWMgQnbs2cuaqT+cu034dmFl9BBb7tMNeV3nsUqx8YMdJfkC0OF9Dz2TgypZ
BUVz8RrzwPHHBa+jxZLipNYGoSUjiUQpEucepWoj8sZyzPOoW4JsH+7iVIYZxhrl6pHiNcw+w61j
jUwMnfUuZKlr25uaVB8uIsnFgbyhtkQsfSSI2sDw5JqCtxtNFtKsEajCEJOoWJ1T/vYpjiWTLzhu
dgdZTYh0SYoU4UlFU95KG3buodvBbRY2oK32lMptOgMU5QkSIHbCt5jX0ph68qiofg/bwDgA2p4T
is3VKMNR81lsRGl9vqNjYIZPCBJjoO71xfgKOlK3rmtVhzBVmuPXedLdK/cEaiEiOQGnr1+IzyH0
yGaLwBiOCFH0VZNyLebHY53LcLO0cU+FF4gaubcPLAW+ckieQo8sg78w1h28lgJxys63xRwV9IZG
dc2aw+54JWwgjhkRGcssJs2sSuymbQ5S8RHQBD40VnmozU6iGLY6vF7o19HsgKjpihf+0W4/x/cl
c/OCQ3Oc3z82J742WPQPMthaRofnpdwPLJyZ4isceXmCcs62b4rgR7Mq6bKrh8RMFiIyu4NWr4mt
VcIzt2hlbaGqUfobeM4lPkcdp6/u6TbCOX0zb58x7s77h3AnMRSrfzEBCGhRxWVgdyFFTLWo6m82
rBYlQLmcpjvgYHJbHYnHcoHAjZWIcszGT2lBPuRk4MwNXzm0dmkwJYp3uCaGMhKgwTiPS87+9am9
NDq7iSJu6z1lw/Ibhi6RVBhcnnOdBEDADaLgx/8a19aLp37n+VwfYwOMi0pIjUdsSdbBm9+F9DNz
yBIghvfOHLkWeMe2yVFPvas4PJypOGp7iEIwUbi9EO8QEAWkD70LMux6qAQomPMzCgMDmQfyl0RU
G7nwWr7Nny0XRvvzkKtA2IquEw4pSgD7k/+TxRDwqiQbLjItgYLbdAsVitnVI/UnyFeR8ilRgFTY
T0wYIqamTitG8713Hzi0k7InrzAv5zdKeSje7AviXR5/AZsGI4vZRyAoEsNxJeRgKq5q4P+0S5pS
7mMc0UN18u7W0axbXpGYMsC2GfZ4/1PfGIc1DCZ/da8VPtrm0yfqNw9qpxOkaXTLd0Gi2tF+tJ6u
xqQ6kkQdXIXTX7XrxchAaJ0FfvHdf3eQEshT5DUO8pSj7bfNfeUdwoPVBV4UyohfVGsJ/t7ifVAy
qloG+i/xf2ydA4SY4dD0KPiJhE+CmIWxDO58hG3HjL79ZSL4AdjcIlBsbkvrePnLBht+rOjIvaXQ
trHzhjFMXIkaHu8ygAk/GF7cuhMuCMOGqTnPMhDCGHlpwJXRB+QBZPaSZWDbnY/H6PMCk2U9itJx
44NPjd+/279XKVMO1MMu7XRG3NDFTEE3w/nZiJProeFXmiilC4Te2iEd5DvF4pQ9y+uixFHIF29Z
THmfhsN5Uf6sNtXRXaMO1cxGzvOT5VridaaP2gH7XgEPi2VF8afNV+T3F5DpCuIdwDTs+SKr1E9e
apDwGjzIJv4+2ds5wL8e0KcTftcDCHkTnHf9yAHhnMxlP9nG9hQfGqYLkIUVvYRDqq25oKxGBBsA
+FIEegjytZQG4UXQQpy0QJWQ6+MlA2kCphg14rIk6va3nzFi44vNEfeQqzu5/qC+j72iP8KKyHE9
/vjMY0G3PZXwWP6LExevewQNbplL1vIaqXPaCCb2bsAqtqVmAGLK38tMSvIPw5FYOzwdV+H3W3Pa
vCJuHco5+R1qz4A4UL3dg5fdozgRFBOntq9zHANeCA6G5LCKF4mvodhuV14xImKKv2yU4oZo0X3y
6GpgLASvSVi/ja4xTWVql21fU2gbyYFdKcXmchM+0uyYu0/eKIuO+duWk5ZTS9RrGc3tCWBbhWi3
b6ygJYVaC93BgPL0WCWX6rMcsicUvxd00+g6dHQ+WgPo/I6E6LdtAXgnDXdZddRZsq5tqym4qab7
qa/Mz5UT/UyPpyLIaMfQpSJPFC9lDWAZ+GRTv3mv+uokaDVaMluG4Vo4Atlzw5rrNePTa3YBEhTP
MNIKhalT+tQQsiSzuJj7fs9fETYs5dLBA99mEbnY70ootwWBaE3vPOvzKqbgA5vy4irN1MMYpDvW
90/aUtPT3i26s1t9r4G/GQKdl/+HKMdgqgaooL2aRKse/kSA7XA89i2D8LPM2gYAhYbmvTAWtqY9
fwX5oo6ZnbXxKbnhn7dMmm2/k+lZkVwjRC9Dw6WHMlswVgAeMszlnOavLBddk/1LnnXR976UVO2I
Ew94gniNVwer7VPPV7yXUQ1xkZzADBntZ7tGuDRk0MwG/Z5I6eHpBTMaJT4gcgg1QdIBNZUisO3C
LEfgC0b9nRvQyoZCdRP7iflgxWiSR+CLeCZ1HzG+MZMNyG2Pm8yO2xbZpYTK/L33w7jD46r0wnKT
uFfyH2J2cQZZeQjGdXAmRVc8vaeH2hpIgHdbCfHELB++kg+qMA0OChRub/qeq28HmF2bOUXEU8Xe
R5ZXCChNC3Bv7/aK5SKqin8hq6kCjLLwLxu+4o/CFTdXJDE6jK+B8CVg0cadZD8z+C7lwQtQ4m8P
yzrYdWP5S6uwtojDUORAn3n0WZ0goxqPYJf3vAzyS93HWN8N76PeMmXQL2rOGenLJLScSOkgeYeE
Qg4+zMeGbfavgko1eJYaTm9m7NAJrqfZwKQI9IFhJ4itm3eEFipr4rhJe1azxI0MjHqyRT2Vq7W+
HmQ5xOGqEcSRkwxh85y0gSPMcJ4wkvyWG7M7xbspa7n3cOFZjmesvwi6yFS/+std1PGWuSesLsud
N7oQdNXsVLN1822IQAALahLjWFw83rvT3aEICqEnTOPoSmu1Jg4Yr7tvluForD4fLs8paL5tY4Zt
N1W2VXNs5DoDUG3vbvm06c09H6hM4Gr50ipKDbSGrVmzfVMgcN+6TAmaiTZa2IU8n7mLgNNPHOa3
Lx8wbSIfnennKmps5ddGohAZq/dSZPsqyLDk5MYH8wwdYiTPkC8CMZO72/1CdD+4TZWwa/h+PTCN
Ckuo+fsTp3aQHy5ydSd+snNsTd4qQ1ze9PMBZ52iJakN3Sgs+Etp0ASR/dfTklXFqEi5vSn24Tin
/G9K8fIXnpJIoufZ9GI+8pd4a8Asn5AG+H93wwMy5YrtiTeiNbXy8+m1CZ/ZljUXV1QrT3+Wbv65
+66j2+Ea1grgJ/vMGbiMSxtYRlRueq6NBmGPMmvLHvMAiiTtAqwZ+7ruH2cBr5XFWR0FFA5cL/YO
LQTppbEIkVP3NUTbg+3sOLM0+rUe94gZVkH/Gqoi17TKU0o7LpE+HEYgQ88BkIf66pLz2i4VpOKT
vccJw+SoloFXWdX+tGdsnDvr/Vuchy2ap6ZwZz/wkx+GKO8LJWLduIMirfUEwQqfO/pMV3JJZyRf
/crgK5DSb6Iw951/momPJqCevNwHMxCXQsXf1Q0P/gFeQZHHCxuEt4Ht5ULvC8pq/KyYn2YMtKpC
m5lFq+frtod9hcUJWESGOkhHfKbELJVFXtZiqCXLRy6pv1LtpumT4Uhv3Ozfc4tD7KzT2Rg/Fba2
V6qQAc4cHm1mv9guNMjyDwTrN8iGoNx26qn42xPivfTIsoxNg7xMDZPLJ0eqVqbyzHCdS9UqHegm
u/Kc3bU+Atl1qDeR0c2yaVRyKWHpbOECjL28ZKephNrkha8jgsyYz3K/qgV8mAb37oTy54yv56cZ
c5spkqmhX4Pu8QgN6V+ghs3zpDGD4NZ6TwNiIbmFyFsYTZ/XBar9fWU6cfPKbTQGolwGTtikSfRV
6bQGFpWGSCMWkmn7s9ysBMVH3wE4n1J7VFA6PETKvsKoBgWD4v4RjvJcpZa2N/pOX0Ez9YPEwvpt
unq6BHZaO5Rj1zF3t+V3dnHiaiHqgD8aQidLXbbTyvIWsR/eV0eMWCcBNoXYgVjupdLQNLDYk8Ez
l5bKRF3MSpB5Gt/Ayd29/yy5rGkxTf7SpuPYZLFC1JTppuV2Covq0Kr/HHqLD3kbT9O4ydoyAoDr
5Gw9x7UIuw4k6vhe8ujePxVnrOf3x5Ybvu2TejiUi8/aGqikt4m5C1l2TqAYtZr4neE31Exd6NG+
I1jkfbzx22dcrRarypwJBTo6+gxFOkYe6IgtUbIJsGxU53dGJcUrl0IZk8lAt/24V1jRX4jSN4Su
HbBNc4iNI3uZqKbMIOzSw+STtJvHPxltu66ZtQ2GEJDmz0LEnjxFszYXq2oPTyeiJr5PnqAFCuqJ
pKSDMyr4dGuv4KKkHp6vUs0MCYKMG62gPMIcMrUuoJZdsmRIog7lLWK7l9iXUef8su5lVV2x5pMy
pO3pRndvI2VV5rewrE95/JMC+7lWA4PEw5ciXUM35Abh3JG3eia0ryIuZsWLE1nJw4d04VSz8WZK
Uxqg1T8V+84ICesKhR4vuVyaVVJpXXD1GgVbYIrmH6umnZPrWOg4n26nQdhdEQujF848l6wlKBA2
OLjtBmZsE1r0zbTAS7azZJMj3UinVNZlbHsvo5fYBg7qBNt+SH4UrluO+LnGLD26QhM2fUEfsieD
4i7/rWFCheP97LBWvAGUr+QawqHEcrp9hd86vo+FPPdezEZLbn5FKBRYii8qkpmlD2xXpFGJSdWd
wDoR0krDkjfPHCrCAjSmWvo56eSzb4d3kJC/JbMrcleaiZXNmDaHdKxlBNMpeb6rzSATgewrzdmz
RA3Mwkmy/pfN97/5bi5nI1VX01RYo7dnaFu/ccKGZomJM5u+xkP9oPkIqMgiNWxefBnnMalFVKeA
HAV5bd74Vr/goJWN4PpYtJh1MakSJjNs5pnhEBfJFNnR4MhApJHT9Miewg0HV/r/LhHStbULp01F
ZJQAo27dX0sOwiSZbPtpJipmy+CR90U/YKi1D42hKd5EAWVQvR/crRaLPng6XF+NEhXxdZ+L4eqL
PRYZwqsD4sPNQavHFrEY5xISXeVV0RpY2z8pKm2J8GMlUeg34ttvUlV1ez+wqKPYDloqh13m53eL
yskTE1Dp2RoC5x6jf7N5gru+wSgRCv4vUL/qnIjEcDGgJSLvU4XVG3hkCrkA430jhAXVhX+DWC1I
Q2sK3h7378hh6Rn2uD3d6KwrVa6jm01vlzh1qr6gbjN0VCygdxvZrIcBqVf/TmCiRnxdiPXgJxTD
lTmsImDWyZYArFyiFt3QWuQV5B5k86yn1ef6mOJIasvTsFHIPGpaUNTRZX/Awjt1QXSP0eL1R6Oq
ni+qhO9uGCSZwieA646m8fdBXiLzHtwRPzi6g2F0yrh0BbIMzkwJouq0v3PPnG+0J/gA1UquTuFG
23BQL17mHO58WdH38m70es3OxbqbEYO7YNELAVRwelKd/hqp6P8MeitpMASk82uf13W9NzNsjltB
xv6/fGKn/nPUMrXGVUTZOrIUioqFjH+1tBrkN71u9i0jnwcD0w9arQzGgrqNxynZaAwamjKzpGFh
GJnWWUy43LCmH8BvjPhNq7/yw9RSdfn216zPalxPBHiQY1ISf0aFgtkL+Pa29BdcWnjlV8+/+FKb
Fo0pfzuriHcLSr57i3mXC9d3sYA/ZNhGU/zhkqcSoqfXM4+8un17kt3HBrSSGj1Iqoy7vRJx71/O
vo1iwnt7jXyIwDZdTR4RRTLzrmFFCniAJeJ4Z4BBLTpsOLI/O7xhuSOksuPlACppSXPNR49zy3JY
CliApYXwv0TyK98GOw/YG1Mr+H2M7cBB1tc/BH/m0EoSQiytDcxUKKDPUBYTztVeQwJdEQhdzjjL
V+th2hVNjT13ZzxFE5azZdf00k9fby6q722Qhirz1DKv/V69653dIE3N1r4DFPbVgO/IMRu3Ufvr
LiNjbu3/3Qi/Z4A9ibvzIahlaDBzN6RiGzAeQpMRnnkud1Ioe9Or++P5l0m5NH5QmWt9RplHnoEh
YMk+KM6aoSJi7iDO5LcCe7stzEwYWP1gy7iU1iJEI9qA+oeSo2GEyB8u5AnuoWt4U20aNW021QC3
E5cfaHv0dmHDt9rcY3QXuWPqu0qzb5X20Fue3HiY6jeIObeOecaYsy5D2X+VPemHQ7SR2oanIF2G
ChMDnOGCw7RykfK8JomeA4Mg6YaDDEsFpy8vJzARL7zOxocGp9jpSR9mtcEYtOIJ0KO2AHmy3GBk
9emRkDsjxikg/33pCtuyJ34Hj2Ya/J5zvUImPAr+t0xneGWZ60bNELlB6/KDk2a0NlHi+/DBxSU2
OftJSQYmuaN5X+45EF/0T0FRlGbw6U6TcgBX9qknzBa/ZaalB2V+KYPP0NVOlhvR4Fh/tcsuRPQU
0O3H9hL3DieJiBalZ5nQzzwsE4mGmP6aw/t9qiGv6EEk0kcvuTuYZ/adEEiQsvOAM7D/fR+EkoHC
4kJ/wyvjaXmBYnZRJXGdlkbFCObzSd0so862RwCtigPDU3mLdWI9ekdpC2MVGZTspDrxqVwiZZAL
f5kl93eFxjblu5XfO8EgETHh4x2XV7qtuVPmsMtNXOZZEZ0q9plLA7oHBTA2eEAybo9xeQdJRJia
1dTxUJICzCFCUj9BDYivSgXPSXYzEv4jjYeAzr1w5/jW8upV1NrQ3vTfwRNIT7/VV9ptSJP7+R5x
omYxw6cAQpOFR9wL3ZKrl716wzogjjsDMXsbfQ649Wfp4/Jiz7+PQYGrPiV0jtsHdJjZ6/R7DnRT
PnH6A2axFtF+IRVDjHXYLCU1zIOekljsoBd35wPU95PH19UJ7dF8Ot9xr8lPntXRhw0hyeJ9iVpQ
C1e2Ocgnai9oK6XWW51nDKpinyJzgnxdia9dDC7HXZNmCMVmgeGwd/wvof7P0BoafEDsDUTNuRtz
y1khsZsm4Z1Tm4K6U20MLmHlGWaaextyp1pRktlFlMC46W8ekerQlosAaSiyD1/LjICSWaKMUoWY
rC+4Vydnu6YZYSG2QrfCu1hEWndyLn9RckMugKUw1G2m56bwlmGP79eP9IrZXWYdz8GD1EBy3/FT
aJNBvVbKkDHhBL7I2wwsW5Bw2UNrLAS7ZvoKRX4ZzKKgL8YzU54b8+fHmzdKO4D1Y+MPqKEGvwy0
Onv6K9NZalYSdZgYwb7OJSzi4js2Wg8kSXOwU+TQfN41QG4Pxnf1NWsMMlCLGNrc0aeFLVDfKX6Y
YwjCHHN86EkYIuu0aWN8U1yTKUBmC/gIqx7FwnfckZjTNUsL0iZvQrtd6JW4BkZz/YmkRLNFvpe3
JmeLAreh+VVjsUAmdmBtenB9cGFAbhnT1azw/Han3qEAPHgCB8Kfv5bTvSeTCpoiL2ULQsikHdBs
y93ytV0SIhgv+zYGYqGZJdHUDUmve+Z8E//LeKZ6TNAcAV29SDFYioKvTytSzx8D+HIkph0NlNtB
i8eOAtdn65cyRF1130Y1ZQUxK512N6utAedilyqiRkH3RVzfzHbsNPL6wwy2j/xKwM77sDuKJNWI
vW1OAk6Z6/5EYnoQbTSCkS5PFq1O5RXsQNtYFTkqu7Fp+TBf7VDNnYn/9VEy1jZdnXZRSMTR6XrV
WZEd+oKmiPRkK3t9pDDjP7Pc5OBkwJdnf2HegbR45TkuPIHMtvOU1lTTYpfpz3tmW+fvKfnR8de+
tR9aPkmwVkBMmWdbmBJDHVWi0qvytIgc4NEjlgO5Q4lioF+hV+epT3XyOSY08+VlU+TXLPGXj0le
DU2ooUdp0ZCjqnAC2qRs3SMl4qQJaG9HF0qkBgeOEjlLaJkNGl4vl0KrseLFyKTNR6i6HWkYzcnL
fK3zQ+ygCcqI2QrBf6CkLD50M2wQ4O58VAmQN7a2jjD5lJJM7aUcPvue2p0f2jvATlwaJWf4cBgT
xt585ftdbxmMTM5hXhWKlZSefr7RiNw/dZgHzPlwUOGPhPlZje/kIqe0YSnk/PXExr86M3gG58ZI
Fhrg+M/xZwcrNv/CwP+1bpXcisgQqmzhwEgfX09RQ/VOENt9b+6+daUtH1pmJy4fpj5tramaQJVq
0w641Grf2RO/r5Rq6BJhIn4nGA+Tiku9aHgiJunseae5LTDWHZFXb2OYPyzPdYeYwq9F+HiduM/e
P0YF89Xc1kT9Zou1N9qtNiR8ztxaZpPY7JBB+kUXN1XGaMQY3nmLUZT+tLWWshZkZ894Ok1gyQG3
XqBlT4YedBV08KaJ74mBQG7uqgJP3desP5WYaeBpVZXY3hOu2snRPZV3goGeSPc8oDVLSj7XGQ94
HuzC4oClFdJ68Z66FleUUSvO3KsIGnm4Vu9tct2Nd2nqsyBPVKlVyWJdBuRrluWxwbjjFFZphnTq
t2Wt5qnvdRjt7xPhmAATIs6yflaDUryV4nYUZ3N0Q2wORVOVSipshHhN32fj7OAeNU/5C/uU+M/4
VQu+nyDIKKO5pkVXBzTXK9lrzptc0/mbIsTGHX8Al9V4jFh4IO4yLCMlRGzHsI6AXZgYXBlV8TGV
ymCY4ofCqJ111KAiwUzYtvraMwsQsUEfyANPHje/bT4sdUE58htM/mzyJxyB1fmulOcSd9bwqs9u
njdANqpvPqQcc+FfTMajfcQoQ2U0/bjaUEIa0H8KT81JiPotdKxqYubRP4AVJB6/4QuWA+fyBKg0
THQNZqOyWKOmAWhIC+hli9MYiZz/Kyjvd2ubQv8l0SA2wvuRntCsVITDbWYsRSyA989HdCn2fgkc
3T9CUZMW4kUSBZWdfGv4rGdW4maoRowyY9858vR4UyGPZS1w9GYFC9q8LiN/MmU2XnW/Spdp8aA8
rn8tkHiEsJZ8NqGxlAxZXFUxRbmVnqx/m+0ZQm5KS62XL5hrcQcSOAPeVU9zKbvwgKejlbSjfwkB
NufrkjO0phtxC+Vlv16C/YUbjqhTeuvxXlhnvtco2NAEsKtoJs6e6ZsouujP9/fbCr5AsDCWd4+L
aAKallDeHIP39yPkLYL0ZjGDig2hQCm09DlSPiSYGmhl/2FocghdjCWukQJGdQhfUrQgx45sGvDf
3rb1NOijc99CJG4yvAPyaY1wo+UCXTQc05JUwj+IKatgx3qZ2b5UJGyGBG+S8WeSMYBshnBlEY3U
fIfr9li1zkvYU0k2l7A+srUDuv/6b6FWq8NRqxkOaHxWzQtkQOILLVAepvq94qWVAJCdRCYp8Z1w
7kcD/QlgTtaEU5GuNO0Riaw/7NZxSGYH3gYYQoFI3e55z9lQOe9WzQNTF1cCkX0/moEHm4BPK7HO
Oe/Pb55V8bHXKjoQwSAJ1naudFaGnW+2/7Z+ow6CZOAD24hdlO8U6bE3y8zZ3fzpnQB7H3pMx0VR
oDomk6PN4ZZoh8xgYIvCLKTW2awKjxZ+o9wf9tHKM/b5+uVaEaAjBTWuwrdd2e3yYhIYmmc+C7Y8
fYGAGU5agKnVZM2Ffjvac4lsIRGPMmMT2fPjAM2MPQsBMLL/9mRtnGjXPervmvC9VgmmJJBdzCin
Gxg+hlYR5VHC1Ft3yM51CGpQjfZ10YQYW/RgHixILAqHy0V/9VqhqfSlhoNBqafsSeaTJyJey6dP
0jD+i5jrwHpqqcPJieQw8kzwEjWPk3ZcwNK5hwp4uaz5Kmy/lLl+MicknMON9n8xMCGuZRP+/KHU
EsGpVFtbLgimhDIN//zbr9CUd5ma8TsRLbODRcBAUySwR9ZvnFAqWDi+2qkw9IPMRxwFnDOtcnOL
7eG9GBEnit1B3HyDlkQpK1/T1OloB1QMYPbEvx3R0kR2d5vr8ovgj43HJdZOFqRoQnmmMTI5fVzo
l1e4LCW3cDpm7wZXtSdg98IoHWhRiwKQUurzOuwEWXMPqpPqhqWL43x3MTEMB57uoBeMMwfdQzyi
cmi2iM5OqY1O626twvuT1KiPpeEWrqEE7VSvP38rE7iXQ8qEiQiHUqnS30f37Itf2ol9w+09hJV0
k8kQCPWDGO3BNBFwi0M2tm1ZXqzaYOYbZuGiC9wWsEG6oiCCigRoEzaV/rBNcypA9TAgigkITwmS
3QXVFZqawSLl/9nEcrbxonxaXTLZDL3eUzicygYUnQRXxHhIM6IumZ+2ZZiF4DGy1Om8J2QQCQcs
yrBh2nrB82+wr/v5qt/hbpJWm3u08WAfJBdWl5B51axkGhNTKAfzPvAEC+cibnwJEhpVRlEzsHZE
BZwQvG2hfM+5/N0CsTEDBh4daLTd/A2dXFAww57XZVSeK6QycvREhOjNUVAwyZnzSM4rI8yyNOLw
LewkvDSyJHFkVKUcm6mp1hfMAxG8f+ZJPBZ3VYwoC/e7kVKBRYofWJqF4FHUUYdgmjzqB1WfbB2X
knoOp2C5xGNvXY11EDL/PK/ktQazGRbLxuwMlMn1cv44Jeo+vOZYArk9PmItFJv/J/Kuwl0eeBID
tLZ/3fmtGbR/ZvM8w2yVQkb06YXwZTJcNzPdgcpkWofHQ/fWZfwM978q+2/b861+H8xaKU8KKQyK
tkuze3wpF3Sck/ajhS+E/lBDdwI3nBnQgGFMw8BqYu+tBxzsYWzTzQY085tk0EvmHnAS0ZH/ydJu
nct+72VRUaI8mZ+Ix6pOYYNslxSJpI/R471T3cLBxihmNmsTsSjnR6kBvSV94nmKrYy05oO7YNBK
LqdJ0WK/0hnngxAVDV3nNX+FMllSfZ68Wy0QDIR5wVYXT0JIjLqXi3fswnLLnDpK00X31cb12CnE
pVja6sDuobf6EfMQxBE41ru9EilIkgTKKrF+OI0v6aldVc71J65vJcRyZATjEoUOhJ2gdwYOWPxt
gK/VXbM7pgOVYnhOPldb0xBTdcdJ5QBX3UN0WZW3gsxolAmY5cJUWY5DnNoCEeQRcXy3DOl8sowg
XWM40HkNJ4WfJP7r/xZm/MNqzCfKVH38AKDsCgiEVj2DaSyYblzgtkPcgJ6wW+aaXo9y5fyJupTG
9f5FgsWP7w4GnSg4a0R3WF5Rf6WoVEk16vYiIj0CCzypL0s25XHqJfrssxurrWFCl6Sj+lAnJeh7
99DC2Zpu69VtdspaaqsdnvVTRb/bP7zpwnoSGRCkHdo3BuxcLU6AKWsKmXwvq5TTOUI9xe2r3JsB
wHYG9gS+hR6NzwNJJEAFtppjsosOHlYc9UgjPti7L6PMgSFHwuf9sPsAm/FWK+tAts+/eGoWOEQm
hkyyTHQC6bqkHf9IQfQWoTi+sO6FOGYGIV8ekf7EEv1EXXrS8uiTSWsFicaMPhniFSm7VuflJeaQ
l00HLNRyfDfmbNa7PhjsBnReAQqm+sXFBnPLhVkP4vH2yCGb36pV8yR3MzNtU3MDhIfOg3ja5xkJ
Sc2sHu/PBj0Z3b+6PiI7xTehtY3HBE55GnHHevo0sl/KKG6yK+ulyJ7KHIKJ5F96ogR+vwdwAqB3
uZdpsLKtcXeRIQysY5Hg7V5NJP5pWdCq8fOi9ZwglLpqd0KAtWr+vkM/TjpmepxTYPIrtG77y4Uz
ISiHJu1OlVZy6QJJQf8y5F2tyocfzLt+ccIdoGMR4PN20Tsy7bzfbfVW4GwFei58Xx87ZI4L0VnB
cWvApxOU1iJg72t/Mvc872Pq/x3igvnNMxU6JCkz1nh4QQM2W3svlpEJRtUelEWxwhniMbtOAKYp
4XeH71gPHDJOLJhx+cUzGXYtTcB3YRw7q0t3caaUqjto/f/samPIHAagIxp3Hxrr3QBBaF9MwILD
HVvyyzfftN023NJ2p/K2IOBGBNkpTXTV0T6f5i8uEvzM4TNIp0MSKZIOa339DX0gyo6hsHatkYfW
XrQCF+7u3nc2qGVKRQ2WWRsZgMJj/B+SlD407rBNsZr1uJx6d5LCsoE425I6mCxlSYUWlWi/Q35P
3gVqTKrP+kCivRrfA8tGdobk+M1BK5UvCjWSOxOlt0/XFbEPEISVC6DvFPvWEzCZNg+GwS5bGph5
j6jmEM12Xdr0cNBOA7fSFV7u6cm3YAlklP2BB/2YV3wdu091RRI780jtBZwAsC9WCEoSGpylmzA1
2pH7stg1juUL0h4HQz27vPJGZ42iCo0lVbJb56DVMt2Yoiz+bLkFC33Qh9EBAvl0C3H45LtxGBoy
3ab1NueREEtXZci+n6JTivKkOJ59Fz/iWh9LyI3L/mH2kfWrgVajHQ4Jg50sBUaS3vSZe0AYegw9
Oac1uZiP0iaryshVSplDaREIuVoENpceK/SBjM/OY2BnVAFjVLmX3WvDhUh1gYYhJcWZiJNU5AJj
ox2YsdRSHS122Vh9szYillOLEzV9LW5ULz5rcP7tGWM+iBaetX1iFVfmxCZJ1BsHGwosHzw3l3We
0IsA4MTtkd9neGGZdvLk4LX1kXl4KsaMVHAbLPZUsw6rERsZAz18CwwbwKJDykiDyCRsEw5Pp77O
aVVyl7YI24DHs84dNgzRlCSBMdANqO2g7oWs9htlgbfdoS6azWnODWRGlWSfOm7TBQeUatm310Kx
pqI1nmJa90Fbg8Vzsko3DSIBS5kP/jfTZj6TgEfLJltks5/vtCmK8WKqH8uf2cWiupPUt/2c6l//
EhMIEXranHH0gUbf1h3hIEXFg1cCDXmd0p8FEH954Inhfl2rdXAMRRaHn+LUmbTquc02ja4KRCrN
Y6qcPTcRcOHQUO5R+e6fFvSKWIJegqoFxnkaGaZfndtZkXwaFRgBDyqZpyBdoS6JlRLpFfP1MS8L
qMrxcCLNiYnHUsb6dHDEy9iTAXXpAAVMWx5tOfy8IRMXF6HcWDQ0ooKP1PQI8pZf9gGIrcd/B4b1
ietj1F67k5HF1p9iTMqzHiyWWQKT+lwDkdS6ZLdW0U9RaBUgKUO0KiJSpOF2uODawEAY1s/hNJK2
NVKyT4T5hulcWPEzduvslQDkjGKkH+Md14RNFRpaGqxJkR+l4sX5Y5U/ekn/LPTIG0kFunjiYXV+
dISYV/FfquICN5y9P/zpchrUZqBYniOaupXUTC/zLKqVxrr47wWd7c5L0d+VRDp7BzzhpIgUq5x1
Uz2SiCnEtEeFYnlpyOdoRz/vyidswG1wrCVqpJWla6BpVrzlS+LZj39UQiqjkMXt71adyaIMmKaH
Nhr+yxizATF4FfKGx3fJwTIbk5/KYF8XvYYEL4bFBNPfEs3skzkhfoKReAvAAKVYBxaQj4ploEEh
heLVYXiuDagd9rNksIXH1WoF0+NsugOKn+8pWheNPaPbg1O2xZEznMJ1olHUW9I2aA7ViDbIuzjC
VbZLQBLXHmgyf/7ucXItNOVqskauB4jBa8ZCFDcKC1IIBNX1GI1eko5rx+sfUbEOoF+3rPCxHdMc
JTiwWCGFZp+1G9PCH1lQc1KyuSllFXq2kh+2PIMziQJj5ohzOh44OdL2mI/hnox/IXh/mNN0uXja
Eib0IybLKenla+hFavUkmSmQBiKR3ThFk0rpIgDrOE0pfdBmtPrQ8qywIQGBd+34NzEG8864geU8
1m8Fjuapk682ngEy5AKyBxYLOK1xjaH5OXn7/IB1rezB9suc65etU3ywkHpVaSXJlep1dXp12bLD
8BI7iP125pYr4KLGLria1AIz/Zg3MRLvF33BNn69/tYAeRSnzc6CSb72I9seXfzE3wzo4EDMVjgN
3viTGgZCaMaJgdI3OlZG+z42MP8jCow4ZFBtIR3iR1fJiJWuwunr6pNsRR5ZIItquEqgplvxAV1E
vAwYtOfgWNManZX1rlDNkTKZmgMLIorrVX/iUre8JX+BixnEiK4arjVInwkCuKAFNmtlmBV1k3JS
JUnC+X6RtT0SMc5g3905IZGEXyiezEQVDxhSVX/YtoOGPcKqEyZu6Lm0oQYwdCRoNE8PX1Pjf8TV
q1qYKBsyoMYdkcTBnq0C/iPnGY9okMKWEhzAumPje4F2JdtoNE4wrLnTNKJIPlhwaNg/k4n8G2Jg
0YCw6U8HhLQO34yz3gpphXXeszADEWtHzI1mqr7BU43dDZ9bnMsSwqouDLyxhTOC2WZIQfw3qeDD
7Yv1TsIut2gmvOqcWU3AjZODKfDrlPsTj/1uYqXtsh8ZTdeazrdQuBBFKWMgw0CNxazmmKB/5N2N
8BiGjON3D5NnCD7NmPv+39A3yC8+Ix6EyEZ2KLiLnTgKOZnKxibaayN3+2eDNEjygjTQPfteDpxL
LlBBMYtzkDmM2Gir5W5c2BPKn0UL5jnbAFW12o9TSFkvNBdcwoPlcZpuPevDzngv0ADETeSQDkLx
f/utVSk5sKIjvlQ2psA1Obiljputtjm5/SZplrEIz7h4V6wpaX+xBjakhrSpE9KH9BDCZmB2Ae/0
LVwgI4TzvOk9YU5hYS4pW3gifk2rAGQ3mwhkHtgZPYaAbn2qeuIoeYb8csw4+L+6Wr0TgN0b002Y
UvvQqvz3L3um7nVNI9T1h0UwHko/rRhxkJ4WDcoHfOZwp8YBUFLugyQFBv7ZxL1+mLHXY9TGPZRa
2XL1Zkh6OCO0FbtKAF+cMHhGafO6Up429sFQkc6a52h53+Nhsn5NdzPOjFAhPUhcfTF47CJqZEcB
my8OPqxQKLNwPenDL8Bj8zQAic5sYT1LoLVwOsYFolJLTh/xHRKVBug7Z0T0vdzQlrZaSjv9ZWAI
8sneUf4UQXnPrRhx23pByMKLUSw7YsFQRWopB4CPSQOWW+zmOXzHAWinFDUOVdwlAX0wsKeYQlcb
RNPLFUZljF4Tof90ePdm5EHMlJFmrxgdAfbe2s+yTN+WqJera6r9aieGX+8XlQRtkxzfu8EqcbjB
PgDAB/yUPq1aQl3MThwOYo//mbuH6hRQVP2nHI+nkpgvGAUWR8auJbP4OFKB9Othm96Vtn6T9FTX
0NvrW8dC25q3CLq6u1hp0IlYc/zhxypMd/zDjDqkPBfAYpD7BqzkTBD3ob9YcZsvt3wf0SljNTtK
RrzVVvOclnXX7rj36qk2X1Ikd9R03o5wNk1tRMlLLy8ziu19hLVS1tz3xGH8nL2t4pAnN+3opvsq
oOuP1f7uflbzwVYYJqn2oG7KnkHT5tVWg/WUJPya5YAGMbnC3Tg+PY0IwvTYO9F5xuVMqFlk3c0p
owobtZIeUaZzrd6ZYVDIRuadS/xNlJuX/ph20P9mOUbpkWv5uVSNuwjFDemyUJKbMTZxS3L3hj87
JsS6E5nVbkNbUlDOfLfgT3LOuQDd3xtX3atiUfT4uIBGZz/opd/eFfR98oXXvSlWqPvKDRUqFz3Y
+4BSaC4f1z5yZGMTKkNAjg4sFVUj+v70ixEDD+o/LH2gESgs3OnldldfNgFqHv3wCtpv+gqNodAC
ogOIKRA6jFvLGtSTDe19m1HuJN+E19M02TZVrxUVmyc/KCcd3/opjXcQBUyb7pVJ7UJ1Fg/gyrqW
2PMNn4IryM1i5ru1TbgA91L60ZLD+wLWZXlCELVoB0U5Xs8aKn51HM8AAbDjRcvQZ8mNKATuqxxQ
XrIJ9+rP7Jxq64Nm/aUJMthUu0FqQpBgGYZCII9dS1rJoq3+ibDKa3aqufMSdxXmOeq6UyDOklNO
2XufCC/5RDlZeSqonxYqw822PiYz93Vpo9pa1AidYwhWIKO7HcNf5iQFHzZo81l1yG8g6TJa6J/T
6X23HDjibMCiznf5ft+FW2jeKjrPoypwg8dX/ct+c+Wk3SKbh/7fSh5sNYuxj+f7ruRivrhv/WZH
EYpG4U3lRUsbV02C2ZJucmUHvR/9vclBfeTJBiAXdzXdnbOEfWiTuoG9gfZ92eAj7WRxTlTfWevW
KFWFz1ZIE5zXAlLDJKzuCJPGLM7OQkm8/oLeNrYEBHwBe8M8fW9K9O1rzaI/umyuehOIpL3ZYpei
Vbz55g93+CHTQ2dA4BgOYLZaJ+CNMNloT21w9QHBGD2zyzm6PuryAAK44rXsIDlsnSDfPq3lG37y
HD/aJ1DQaSKi6mMt9J/sRTyo2IOSdlGyIlDiDSUh3+VGA1LnDA4AHx09RL7+eivGbSXtuwKc07GH
1cYbbVyy9lGlKY1fHrZ+ANNwYDq3cHkYuMy8eI+4hGwI77OVa4NeGXEhF+xWLOcCddz56dFgkNJ7
fBcdn2ApYHB/d61ZgNn6Hohz1LMKX1fh80y3VEFjGJ5wj/m27aVemKLeUGAaXjH9YQORh/ToUUac
1XqOPLLmcgO4D7I8bC2st6LM3WnlYi2vtU3vtwE33mwYMVPUg55kPDpir6eNZdbXk8Xkt2s+oQC9
itMrzrXv2l8GMRjCTsRVm+KqxGDRMcC2AZO/yO2CYZzBhkmsJDv28G37Hc6ThIggLiEGxsF83BzQ
9JdY5r78ZNfWN1/EttnSRsg1QOQ4XLCJPL2He9nXwVE/4IoSzkhiZTJJa3MDU8NUVBL9isdIRn54
N8dRJtjUsCklhe+x+wQlA23mbDXAZyPpaXxUfYHSZ7vV52WZAlgwP8d2l3p7BtE0NVqQwYanTkif
gf8dn4JThcxTxIimcht8jGi5G1wFMKKG/dJmIlwPtKJ/I9MDiFbiKRbBZrEdjs54joWDkDlYJk2j
06P6MpscCC3HORjFM88Lrhs3YtXc2F2oqQMZ5Rm84UceL3WRN0X0por0BwUDc3bE7rfak8X5w0fm
mH+l0KnCLjL0iM4G4kSkZksr74rM4cCnKrsR0z8OUG4FkabylrrT7Hgo488Ab78uZJt7T1+bs+l2
1UVV5XbKcF60f6ObnZN8ckPz75Eh/gJhX0UXx0no8LRWz55EWHNTLCFHhdTo+S66hr6qLaE65bpR
kAzenWuArHMtgIquBB7y+PJJ2Dgwy184718HEn7OA11fzq/b53kPup1Lt/Yt1QOUxf8McN82UvlK
vCadOdNiN4hIDGsPw3r71wWP9tC2LzNAa39/hU5Z4K/S+RyLx/GRooxYpuhQ2pJz2jy1WXmmq3q7
8/i1p47vCVgzka8f2lEp2UCq7msBOfk6RXyh0y3Zew3d9ImRd0s752S69OfcOkkFGp9S+TTk4fsv
gPPWXB1FMMdTUvOBCyQoS0adfETTxgl7TmgMdKz+h6sNnkFYSvJ88OTXYopcdPAKzTIYSg1P9EAX
jJqr1CzQ0Qz8Q/LvUc55dpdQI4JZuF4lKFRhg9r73GuttNjtewrZ/OITDpsir+9tukgtGowtRkwi
EYyKu5ErMzmq30w0+D+aG9RvrEyjTGrMzJJwKOAOe6FsQwauCyzxbDTNiXaT4ginm6Vb2oWjWP8z
mkh8c+lcLVv3/PAcjQkJ6TfIIDkfNsISO8qRLTMNV2ySmUqt1YSKu8NEbpWpiwYuYxz3nqlyQOkf
acv8wcWIQBmkFJBhtrxIfCnnrJncdfCqWVcN3RxgEiujK9Bd7XkpTogjQw6UjJPZvUbif7dBIPOL
Rz9ouP7lCkm9IIPJiSaQOH3pLHfHLu6JFvy0Sozt3y9HKnpk3myau6QLi+CqRLpL1lx93XNPBsCZ
zI61LyoNvhE0zSsarnLJgy/431OnxWBl4MS2fBo/6odRkRiHspDckOP+B8dodbLp8wQsH7iJs9qB
ClL7KW4GqDVxpb+Ykc7neB3BNm3UnYmyFgTI8PHkdwSi3EqYJ/GhRA7ZLVWXSK+kuSKkvYNt0g5k
Ke0Kyaw3W4iWBPFzelLp1zQf+5etUjXtw503R58oEN0RN79zRRkXu2bY9m6jKB0doGkv2caijyik
/TcFKbmYBfnOZMD9HqTh/zw14PfCL0exbI4PuMmJq/racQHAfAtjVqsPoe4fKAGZzZ51tO9fVrD5
yBTHhW1nGc9NGvyU/H9A9xHMPwHYyhsXKPsZsNWD6Qh92qYdpqKQcb/sTNQAKQcV1xXyVJhn0K06
L0vtkpXx5Ryf0Lv9EYysv2drKat8YsHYr9mm3+jETINVncP5Uou1oFlia2/QSf1UoOsTVGwwSCie
YPDg+2R+bdxLBeIZagKvQzXb2IvLNnZwxYlCFWohtjXGdoob5hxkX4wcx3JxcpjpErnyRo0pwHJY
b554T9zvWydNveRAsD1qyNtQOqYz8yvaksRZf57dBoK5absaf+VQGa538Tp/4q0wE07e+e9VhZFx
LrniTcrHkkbRioCgPLSItL1YaQGr07uiieASTEJk5/foa4JnALaiCtSSagnU7BAhGPnLC9Tcgkbu
UCrnwVDyRgYlDm3SzO/0i+DDSFqvcjipgi2nfzXcFrA03vX1ZX0Hsf/tBk3fRlHOy2RuaS8S2Im9
BiusfmJDQQlLR9OffQhsVFS+GD5LD5GnZMC8OEmjYis1IJWZHHIl8p6dMG5FThZrkcV4YldTSLzk
vm6/XubCCRyLzOWeviJSn6Szw4hy6DUtezNaJBMmELL8PJHwxoeAFcdzYjTNTkkcymdDUGmDQMsX
e6os8m951xvGALSEjWLBVAF4AKbqwLSQWTGzDEBOCe0VrnGWwiHUiClFq7CfbrNDct6NN/oIeR7s
3KaWfZU5vS744JAPG4mvozoW99SUH0nhSrSi0WRuv/1ATRWyLhM5Ni0F12+xT1s861XAkysAfv1o
/MtiGN2jm3oJKQ01ApEQ7uZ1VDmNfA2PuuFmFNgkiz0W7HjnaWTCPZ5jwttLd7guYxLghzlENz6d
bf8iAb14YuszDBNXWC450Fvs019BgISMl+d13WzLmIgDOBWmDRqq3X3RrdyJhEpmz5kYfJFBnadD
NSscDw951XRkZI1oQ6mJVD7PaDeXLMUxbe0wPTELj0zvg5N43NNgX7AzKnryz3C/3JmeG7nKF/tX
JgVggkwdF6wlATR1LDq1ScHNIJQGYyjCy2btYX+EO5CNPj9GA9WkltZatOyrH6bIKDiZjJcJObO0
QK+kzxhPLGUFP4n7tgpyhlEgDVVpjoFc6bO4j+aZzjFPKQs8eEj6Ad24uMFqLwgtf7d/Xpzg/Vy6
YME2VXfVyJ6WJ6/TdibdOUIy0L+g/uCOE77MsKZNJPJEhE+LcPRRxkcJwZ8E809+L9zVxbkIi3P6
8QrzE0ZW7LKLR2cZi5+xMubgVHVMUu327tg8a1uBiorsBpbAjTi2oXfq7yxCOjrN2NvnsCS26up/
hZHqivmJTiVi13ZcCTz4S+die+6epj4zqW8Jmig00sDsK+1W+zvCKIo8ksXM4MK8oPoLqjYP7tBC
yaaO40RdewyKQlqhpZ9UB5yyP1yG5SjKE6KQx3VOwBU7htEE1rt7JMqrPwb11WPVw3Bj/z6A87CA
OUbZcEPfFLzHei1XLWZgLkF5yV6a6DT3Xi5pwdcm3bC0wpJARZA1YEOtIE3QDmWli5pb0RuesOVj
bzSQJNMtAgwJiisZAmwiTpOPVfuYRMi6oPgtpqZdVi/yklEPZRpuDGeIDL8yew7tjuz9vyWgH9a4
sgl7BrQQqhtiP49IdGEQ72Fn1SGZlpXm+f861cQ6ctfb42xy/c+z3LbYTOIcaaAstpy+5hXtZAIp
0JF54sF4Z8+jHjQNONLHelSNybWlTUukR29p8UDueb5EQ9RrwT9SkbcyfCoZntAguj1iaF3W89Ll
2apcb+yvm/iPrT3SkzihG4GuGvKZwvahWO0wgwW5pF/CZtF64xdOGL/jdyIIJ28OqwAqIRk4nYi0
GLOP3gR4fzmXGIv7P6e4a0w7xCC1FZipsOQyld0AownSsEklxU0tHt+3Vd/3TkJf0LXTJedauAv4
zJSLCdHcs0V7aMPD08VXHTTsl9vOwfQTIx0/T3By6IYNKTooKDXz3Nn2ttj9j/Wlu1jdCVZt7oc2
fJB2T1I7244kj+xCN1gPGhH9bZI11vBd9R96ec7MF4ZTqCz2K4ndpOMcovPQwBXXlOeyd+RMmtzL
xZJ2STetfMKO+wKboH9O3kN5XrqVfVI1ec/WwZx2tRlTLJSKAXUVkCtq+YRAym1+lLP6vEEdHrvd
cHsiF3jnI6XE7RnzF3fEDvrDWIuPwbQ3xeLzMFgp0TyhNZm0xKvgTcC2LkbSnmVmgkm+4Z6r0nnY
QsjivxLE2Y1hdE/nwFWxL3A1mEOK7DYfSpdiAijhnzgFZjQecIbslYRImE1m8UZTQrr/C7Yr1zqi
Rd0IRWLwXiHEOi/+WcLBT8ixsc9EK7hIGbRCRHxyHd2USglVvRpG4MrRQDqoxDwPq/ExtTO0eHmN
jymKOuT8v+30PrM4S1Oj/bKrCgZBUGyd9JrieiwcUL7XGAVwmln2eDXurDIAN+Pn01yZn7vikD7c
yMCUjwtpuRfg3lGpOmXCK40znQnzRil+Q4bbVQur7CZhccmAlh6mf68tGUpw9t8QiOAlYyu+NYT7
d7gOVClnzqR5b0yW3fE8mf04Gbj0n26tDIQSZx3CjoX/xW2ffEvCxVho6S62kT67JmaQXoysoyvW
h3IVzriDtZ3bgRXQiOYNMAUNL7cuoybVdwQZ1FvDgEE4sRtuGX7zN0KJGu+9Y84T/gyAPZLBjroe
VxLSs/5VGt8W5q4AQrYNqagLTxZtiyzyp0rY/TtRpkoAmBoh71r//NUyFSrwThNdXsYO81Ks1TLi
a3iVil4x7OMCQ3Q3Nff1UfJLTZpIsoJwvt+NoxMVFo9GcyVDjnPNdWpZCHdInRHZSqtsi7/+pG27
SsNeRm3jCmJ7v3GwN+CWolbxXWUDzOxnMlVMsPXNy6wTPquPYnLNSu615acizcKBQjDAN4LhTHn0
i9PAb4qWCrfnQB/5NtJ/lAyE3R8sFUwfXiZyJoHla3mdVEpCG12owLFQwu+zhKnSok41EX9vpDFB
/9CPfCJZjbEZu34rfkGZZcG53htwo692kayWymXEjNjJnmE2bdOOlPfg+0ZgZdsXFmS7RQVBM4BQ
7V98rreWuN0ffxnnrZY9ps6J8aL8aIoWSBNiRgCFf4PhqMHtIDk/055wwV0bVyF+hChNc5TjIca0
4GxzoRPE7amXUY99Lj6aGjd4geiAZ3Z9h7IXE0MbOZq70ohpIifbDMWRrFSZxAxMilYqbqfdv/Jl
yc5EOrzyKYtBBkztnSscqiq3fs6ox4vPHT32t1jrHocmgnQHddGAR1CUARhtUD7DflQJr1PZMw6m
Gymkhl+5eHeoTxmVtDajTEgZ3H9mWU7tF3md9QJusrb5XIV8FtwMrrCAaOUNF9VlSMgI3cuZ/vpo
v5cVDH+ggSHXANWEQ/ZdrA4d12RaW77UPrOSj7lP1olLGcokXDWUz3JNSKb/iuyjAEawYaALoVyF
l3JpVBimyEYIuvToogb0RNmsYgdgIzhpXOTFzXEfhuL4t0I4OSf6cNnF9EodD5NjNSgQmOGxzNlE
fJoNkz2bGDk3jtHvd4RWTH/YTOagQXg6MqTTaVPT123i7f/Jm0vdW/2me2xd6b2Zicg0bRxLWIkH
PEiXQ9i3ed5HU24etDDb9aBcAMy1WTPsqmnMZJsNr6U0fyhR2aR9Jj7XgnI2DWNTq/r0wa31K46a
9nICkPniGk1cU1kY+18Il3NVARWbmW+TAJuVaTJXt+jtQDQcMs57/lSEH5HKcxe8wZplmCWNsAOq
frEOH7IFmGDztS9qTk9uDBEQ05pBRorSRVn2abanllCX253DHkanBkJgJQpxPBFBWzVrZOVvAfXZ
g7FileT44NqisXEMhbtbyFt2RhobHyxxcQnjbg71PeBJT0XTCl9gYvqwbvUULhJAU9heFYAxTEPu
BimQtpUHAH7YxNSfBa6EX8OkVgTcVujHWFsdI/PRiqCGzJDZt0iK8aNXkWHtwDOjhR/3fhFsuSt1
R7oa+HstiZ8UDoIHvGb0cEcwidjCGWQuRvJ4wAWs6p+Jg/C9fK8tK5nfLSsttuZoawMTQ/Eo0gAe
PRS4rdfftq/37cWxlGv21mHlWya1OjLJk4a12J8yZkXnY4X/ZxefBjqwicOhY+QhVwdzz7F7UgZt
P/W5WrguV5g02xsKdDlEzzwr+6UYjdvcpXB+XxshZjhImeKWLKWlGRy4Pdwqj1olVVr54egQO0gU
URKBvc1ykP0ToFIMncAOzVV7EI+9kEMBfgIC19+VVenoeJT5mbXPQCmghwW3zlT07KbciPRfy2dy
qsLGvM7FZHe7xplyGurmQk/LKWZnJMNTqBEX0PjSk3qcmINck0TR+7IHTw2ifIu4H3SjU1k/wpsg
E5f7OjgbDVUlJQIjnm4Xp8QO7TTxEQObNUijl46Iuv+ZRQH9knivx8FuSimKd/3oQGE5pVCO47Y8
tbntTnhCqQY3MHcsIFrTJNJLraP7//fFplL8PQENKdOWBcdC4LDgqls9kFbRsG26p8DWppui/aHu
+Dzwz4stRbfcY/v0NViY/DHb/zF5fLG8DbRgRmd/3B1bGArEOvYFjGhx5VnzWSBh6s6y9e8VWp/w
qrCMnZOAtMfwfeZJrXe0fAgT9mmMIgfb3QmchvI4jK4lHe5eCaQTxBNlH0kxXlgvLSC6g/FIFqCm
5md2GtSkPFcnqYiQWe6MgwdVUN7icoITA0dWb/I8cohsiWZ/H2nfQcPAqBU4pNUoN/s1J3hRddXu
SX7c9ULKc6eTQR5c38DRZWPwMP5uS06aYm8naIpxUXajiZZRdJDe8tadBNqraKTZY4JooAyttQea
qExfYW4LSoeASACmETkajMsy/w/FAX/hj3E5eSLG0GmCCG4T9G/XBwtvXKE4r/l50qxM50G1sWEU
RUlPRB4m+ino1/2WGH3Hofk8HEZVwbQzrkqM+ZNxQQSI5VYeGLaa4OFFfozX/O7hVC5Lfnjjtkg7
RhLBjg512QhUc/mlxgxOaP4NDvuVInkh/sDGj2368k8q1TM8iV2432JaTTMhT5CFmzPCsD9N/LqB
KfPYFR9ha8JjrI1p2lC5p+m447vMWuYJjWKhM2jsZSgf78tVj+qyfK4CohbTJ9g6tTEvgX+THHeD
qg3EIT/jtZnxzxeOXKePLYDhpJ5gcjHQG/I/C58gnDPlnqTsiLwh8DCK7ZUsigbdW8U8bK80MvPf
JBxx2P/41RLyeFAqVHZXk+LEzh2ufKg77yMZ1wjU0Y0yGHlIeCMCeUMOwax4BYi0yrxNnsaKGBOJ
JIq3+q2znar5yTm2g8c451hEYM7LEsao8EH1pSmWCYyBs9DY1s6cQQ2zNl9DT7MjjBE+S3b0xZqX
vugsOQMpGC1MDMUyzIwxRWmVKg6D7SqtiDSBEmzYy05dAKc/PUOLEgw+R5vhYWrLKMebIbnCwVo+
8QgELPSy6wlJdsS33IYYy1+hRSVRAl8achtrnJnpkEol2EHtogBJQ8MOHFpruKRYUY2uX/ZtTiLW
LsYi7q+z+BtlxLF6PgI1PagF4gvNYoGZD5ZB7XvK/E9n8XgSg7M4La69YpzRX/Sh07d3krFFjqIB
L3l818tsycN4csZX8fdSr4mVmoVuQX1N9FzWAVZsl6p5tLRSzU4x6PioxXkJ8Cyf7X+QurrsdArM
G2W/ujCMvKZIGHjVx0+so9swrHBH5LUC0USrBBUYTPm+9HyPD4WPJGfxTmCt+bpSrq2Noe2Ui/Ej
1VHoKdPTma810MjdG9RqyIszb8mPRbXPtW6+RAVJiUaF42RovEQIHNG1Qq3vqmLG73R6VVeId6x3
Uk2CY3S7UCOOcD0P8rz9+XZnpfE6LjdTj0eEd2BdoSOo7ZwG8bvqOchcg1qA/jeEekVVTWdfNM+9
iNIY5bnT5WVGNIZVkXMg7UYfIKOm2+uD+pVbu5VVMsVH5cIjtNecUem8740O5zNrY4mqI3K+/8cc
wjwSaMPxxf7RiAsYoZ2/zEZBTWTOTMprkb/NSKRlVXN+5qk3H5RCZKKa2BkUs1FHjxX0Kwm17foE
BLb1pprzHJRGJz57uGg71/IFgoSE4r9i7t7WLFrkWkPUgnfpP+0NZQAuZLIXN++NtqwTP0H0Suwe
z8beT94TqvUb1xoj1+jHBMJzkmhoaFsUk00AWFCbVSmSb+3bgLHXUqBCtAFMgOnJnJqF5aZCN25Q
Tp12yk5Zf1sPzCUj0+0jQjDSL+A7Yzsd9R86weTKChGuCv3flqUBdw+olvSiGbM4W3vTbEr/QQEU
bJDyYLNF5uNhNaRPhU8XwLzgV0ec1p9BH9AxtrL73jUCAJZbXSnejg1lhL+TtoUJ/fBV0N2+GZjM
wV40OhEE6Eu9VmJBkF/fU9UktHlQ6fD6SahWs0FS8gZmC1dMfRSaIzEAhp+gHjzYYi67bscqWUl0
uPcYc97CtPArworj7Z2X8fc02f18qFVW9Iio05pJxL3xdMwgKID0yTmljBIMoNJsmZZzNn93lKXK
J2JRFQa7a3Gk3DBK+WtnUjRdoL6D1xn9HMlkm3fDNbUt6t7g1Lt+fEtXFPfjtxAllJYuTwFejEak
1Kv3/FzSy1OV31/5Xc/xF5CbG5FE8JIjaoP/xb6c/Kct5rzRxviddpju9qiNaLV6bsrOV4UeYo9A
0zrYe6flYRt4p9D0Q0N0fD9ODR86EKOoN0LTtPv6gXjBi64hWjXAT7gjiNkkpYiQ/oZlOQSaqvcP
oNLncQvnMCN8ADJ00UyIL7A0KTRNDnWOpV3J3dkiFzWKRwvHSHGRuiTN1AfM/dWheWn/jQSwOk3V
3ejCgMSrYL7WOAKuc7qXw/R5vVRbpTLZq0ZUROOKsKDdFaThOybQKFyLP2hYU7sS+KdXsBKA4u/1
c/qBAJ8r1AuHT/gSq0Xaz9sVKktPtUbxPXZqsYEokxd9VeuJRfR5PTbBSCskcpTkyPdCZv4674h2
vzjqzSkgL487snYcVNu2YZzY/cQLyJNQjaM8Vcff+pWpu9ztDrT6TwmwcWvzuc3auZdnVhtF99kt
8nAhVTLdlhNg7Hrk4TItG+9smc4ZIPaZ5vvJ9Ueo0C1I2rx5W+NNEBKwbvybBFjtYn843kdtk3D6
ZMlB+igDyvsXwAmhEfLSSqxLYwPT3Z6XyR3Z7wUBH1FMW8WxkPBb0RQqGyX6wkjjNb5J4GU3xnuP
X/dqSoQGOu9CoDXIfZsIzLPDMoGzcOToz6UUaH97jF9Zf3Nfz+qRnfk7pZ64ZbucqK9wDzpcA2C/
wUQt1KMAHhw2fW/kq3YKjM0AcJDrohQO3v6feBUh7oUywUqfGqVJ2+ZKOA97T936zKLclM4lYZVR
EQLKlXpvlowxouI4KYXlxjeAYv2pTqLSoNdd4WntOgV//um/ZWTCAdhZupxPPPShTyXS3/N6goWL
cyMPr7eWmwSgKLmcmMkota1N68uCg8OB4uE4X1Mt11NtbGxepivBIvyaHf11CNbZQv4Xa1PLuAfu
jM3c0+wy32HjSQNXsJ8KKEEs7EbYl9kV3p1MGhxUzMS9wXqnFmi0ldN2BH52PSWEcjYEi7QDdj/f
OT4h1btKcUBVrX5drQXreb12u5QbNb2/BjIPfEHrzB4+AkuxXpi5k3UNcgK3oNhFQsukTPNIRk5N
x0cGhujp4W/Qpqa0WOc6PRX+QmrhZGmDHgZqZFrHfDdLZgrqx5OHwALuQuTmVvJQZU8jGHTrFzGA
5cldU3uDRt47va8iEuCdsx4rcYPPiHQILXYK/6O66Q44UUN9R6Eze0WqjSlsJ5r7Yaegur92xkTu
lZSLNQBsShS0vQakdbHdLXIpvt04ckWa/3KnDuR5etVEcoFTFH5QlKt63kMuo9dvYEFd2hDP3geq
sDI2inbVxhfgZBa27MpzeeAFWdDC35VR+kgeNnsiYuwDUakZdUe95JkPe4IculoukEYyXvI0v/8P
ZxuPTXYw6+wsxJcA1RE3fmUPnfPAGPjlVX3Zo+oGq1wa+4e87nTYHdStWR0XeNHlxAoQ2vErceaZ
/OK92hxcorQmzByiomr2AucfPo+wmjZN/3pvQaw0ghIFxvcB4SUFb8ECSUt42qYbFYFVdhegLqd4
gzSaf8bcI6tpdMUQRsQF2UjTSjcmXFplp/KlzyAiGbdNf+SsbA811rb/HpjCsHwS0S74SGCDmV8T
Wrp3wfD4rljVbXchT5IsU+KM6vdrgNh8blwl3ChveyvjfEFXIeyvFuW6UgJmRXqCTXbGT1jzg4gh
/sNd5sgPTO2nvlr4W9ZVyBjav4OCdgspMrHoJfCNGw+Vbr3X6XYxMKTugGfKK2Ta4/lEFVDmqub6
RFfK35VHftCYUw8yRY1zxjzRJ5g1rWjVy801ZUYBAOTQguy413hOus63UULtI7D+Fw3/XDhxyjOB
6z6HM53OKHu26eaJ3RScmP0sOQmpMxTw+LO2vtdap9firyRsxishjzyXEbeu/IoRjbZFKG9XGAbn
lF795DBUrlXNJ3luWH3JM0nsABsk5jOCFFP9xenl+Pvv2eYYZJZURJwrqx5lEAOINWptBeetBSPM
dQthGg8m9uEDlxNbd2qwgNT0Ocwak3EW+u9Q17PikCQGQmy1TEEIlz6l6Sn7dBNyeoHGtv7sxMsA
ZNFHXCJdx6YLP+1eDw4pyCcS3c6LdqYGRYvuOKpX4ULPIMtdYT9gCJ1ktcePeAkSFPDdIcV4DVJM
5qgdHLRbLjhcjlK0pHRY1stLLhDGON8n16XwmnLgvdB0RF5t1ot0KEtYt8wifpisYq6Jdveg4kDO
085I2ctpfE/6ycIFrTB6opME6fiW/5f/7a+z/nyojm8V+AG1RyE6fII5ZAOLNKEwhetOIly7uBt0
23W57Bb0sdZktPGZPL9Rx/HHxMozacBMgQCpmpesR4/wT4UMbzoHMpJ+zANGSINcf3AHqu+0znaD
Ud2pYqlMBl9uQ/gli0rTsnSUMEj3T8HgrdD+9WIoYBPISScwKoERI9fExlXOkImeD9iDmAXExpuY
lzE75MExLvpLcCU1SvFStfAYCKgpeAeXMi2N6TtOr3ZT3fBXhOCG7apk2tfDlXipNXzCr7Pa0LLs
n/9kTM6YS02K1GeiEh6zBBBqg1zP6vy1KFGQpX/atLxh++L59ysqPdYiplmWETMl4HbWZGpr56/D
2ZLSrgtlXHTOHgTP+GHapPFCNmLID9R0aDZgds4GtJudMZvb3Ph2y0hWDA2uqxmJA8b/2gwgVXO/
TgZbzkQkvfzFLCxN0cDHUk3e2ijOOM2BiIqYOkIclu0lsvLzNsytjxV5DR5aeypoc6Uc5CuT23ZU
H4Hm5tfgI5uIvhTfq//SNokcL/Q7b7mmFxkfcVSDq755GPdorVEZPC1L9JORPY6co0mHJ4EusyRT
hJ5atcQEGvaVynWug9hgNeBBIPAwXgM65GhSeSYPOItFTLDi0XC4gXRX2Sjumb0BrpbSJ0a1Ykii
yWcpItuhjbPT8MOyGeAIUIjeR5QiXqRMTqC8QFBKnJEsyQ1Sum5Wl7EIIBwULrFpYq0kKyrWL1Ik
j/5H7gFbgk5SoVkkwprJNuHoYTJ0jlxtv+Qxbi9AGQBwolzoIrO0L1WcgJBQHH6jdSRw++TQPTb1
vqWkyMTWdWi7J0EPBXuAP+HM8p/UYv2NVbWDnn6W8NmC6BxQFwMyQfm34pqcezUkMZeVmXLOR3/V
eAlBfk6AU1yU6qQoYVEupLW3VgLqKl7uniDThcH2fwuMiDauuO2Zoo0jNCNUpktQAb3Vaeeak73A
6vGzmzIgvwIlnx7aP9jx+aOjnm5sCg4byuUTaQSw8cPSwInynu4EC3DABGFgPFvaCDVfMwyLzy8s
EH0K8hNZzM1ny8FhqKuaVLqgEqWUPjIW+PNldKaFQEruK4sFUrD+K+GuR85QvEbvrp0warrxYWjF
hLrGkDM/EqnxxGyVepkPSZolVCDKda3VGePpIkDs9t9kIrdtIOewvBclHbjCy4zuUFS8uH21rMUh
zCOAicxtqEOnnx3TM3YBHvQv9GCfyfcePaDyZa+JwaTP3GJU+QNg4WfbRJ1wDbF1VElYVKkzoykh
AMPpj9tdyIb7muR3ivY8OwcXqmYcApJeM9aeOYrf+o0vukjeAO7+UDQ+LW1t1wfjs8hpXGVbOAKB
7Lf9ushZmGMf/WKVs/mvwlwmP+sNPamX2x8tI+2WH8IjAiyA/zCkA9/+XbJlS0O8Crfjx8Wresd5
0cGValOGu54EXk/+iVi4C3sL/Zgu/BuywfK06+hZo4OgwUGJADyDqnKPp4O/luRYOG85DD5TgVmu
pde3IGGCWKEDTQ+36EEpqjs/sn+3yt6z29T0GAS8Nhix+xi1Xn3Pnqt5CVnPNqM9TNDjUiNKPnNB
lzQeWTnTbi/RspGeaC9IuNMZleB/d+XBpj9yDMBEbPKmNMYx9zENHisiflt6CFrgO8yk1ZGDOQhP
kKww2DPeWT1Ee+Q1N6wRZhm0JXafyPDJzO+zLyzKGOFozijVC+3XsgRn+45hjV7VYDtXKO6LTOSA
z1g6WDl4dFunEaufRE/7I8qcivi2kf+ulm5Hq+zmK3NqbgDMYp/RdTaHf53BCA/UUJ+iZaLBH763
Dd7CeuETY5Nc/Lb0iSSNKNba5Qf0cRGHvFKt+g8RjSNumypK6VdD9ExXp42MrYrYCRGU+7/jdiHC
hzHBqICf/OWTz1PRsj5yc9pJlFL6Z2cRFg6Trc4NFoau8+33MiTi25+8wy1YmyNoI5IbcwyRNcja
F8PlteaLOkgEwJ8COK7Hwj9bNU+zpoN44oFijQIpuzxr2YpveLtFRXqFZ0fcfVu6u/Ld9xFH5blD
CQex6xq9w818DztrlwRYEthaVS4JY0Fx2Y9ytfznfSeVkJe5uWnraO2wJOViBlFo9+PYFk7kWqEH
B1tHvGeLndOeqXtS4ixR1I6gZjRagxVNmj/1Q80kDz1+1LIcWwYpS7Ezk4PaUocapCMS1E/yOejb
bziam/iDwBylNPiiRU9erEXafghSrxd3XCfVRF4SGb+g9m26m/rzXFlIdsSjwRMGK623ni9EIaDY
Tyl1RrzQXYQOW2QyZZSB052pHOmEwDzPRhTIC4iEHAVoyDK62gaEHC2EEKMILpiX6GayTDbUtB1W
0Kb+Vj4R63YL0oRRtv3E9uhmbbYBQ2y/ucrSltyC8rw9MqoQZix+BhMKEmSk9XyN0ZuowuPYkso0
XqvFIb/qFZCYoJ/RgYrpqbZWQ2Rz2Fk7gj2H5PBVV1jn7G8VhvBJGjQyCEN+eVbRWgdMvyrXfd5K
HZvHasOTYJfcjp5y0vLLuTVvTyrHPeptfDrEMGPLIePkJQrTEjkPPscPw0mEUblR+VGaeWjkqwmx
HQXyB8Dwxy0Mqez2z2We29VFrxGlpnnP2gu7y9SQr0CE6Sd5Rx/Q0edFS/u00Sx/81HuHjjrQNES
6sGNDD2k7GQC45Tda1cy0oFeQbizrXf5NCOEYrdXodFS8PYuohzAWEBErMvPi6a/WM3dEMzQ9Gws
1azS6jv3y5426tNMOJsnZAWF9M5Ci5LyFGvs+vcuihFr4d9IPdyJ60HuTWTRajE7UCpn4RbUqV1W
5P1SBGXEFZwRuHhLFOU6EoEHVuJFE6ZUXvDqgvahgA130ybUeyCzDj6RZOhhKiiGpXi5f6AP05bF
fWdaF4E6+0MkFQKmogpjJss8hQNYVz7VkvuDJQVyisEMiQuDjK/9WH6KRzKJCOQOS8x3N6H2rX+w
Xh+Ec97cA+tpTbQtHArVC0591dXo5mrLUXJT4rTnrTg0LgfHBmge/0C/M8hinMlKSfJHDL6IeCZc
v90V4LnLE7MoAvRI8nlLLB1UQ2jqE4SOGSIhPkBFxlonozhEhrzLKvVrRJxjyXim62NHuDDDuoUB
htp55zl+/3UhpY3+7T/bK7DT6SpEZhmMX5RXHEq4yXSZK4d7a6zYpTvdclNijsaHXFZC0jkmDBWe
6rXJmQ7IuM4pmWt2MY+nrhjX6RL2WZdb2jtCi8XUqEjqwBjFa+wUs3wW9pUHbON2CkEGyFp+MwrD
pczqCdUDlxznAyH7cQJVF9WB33WYcEkdCaE7ye5hehwMl26aBXUwghQfUo2Pp4S+c9L+BTfZJp8R
oq6X1ymRQbkFw14rsfTcLqsC0DpPpnHCYf5rwbNmgDJkBlm1TJe14OmCvefU65Qv17R66ot7RBf/
+aGelYNp+n7Ie0HcYlwKbDykJYHMdzWytpKWgxmdAyQjDlLpVr+W1oBUl3HKzbbbXTy99CFoyUpJ
b4DelWSi06PDqiLwIIgVUSjuqYnkAAuDX7QTSkSEiLCcY9w/V7fwxb//TAUnZuSHmOE2JaWh+sNu
JB0zHKVORQ+oZRYkKvGKZKHtL8P26ubiRNNrHUo4raD35bpNBfoLWQNsFBy3J/72Qrb1KVGAt+2q
uwh/UkqTTe4mxjGsXkLN1TUe4s9LoXusXPFOu2euzFMdoBHwTGHu9jV0gOrH34U36nnerdNGxtPW
GTIHERza9FPBvOw8ZSGFF7S8CGMWL0p3KaNwmBFtCjO+gzJQbpC+GCeXvxv8q36t05u3dI+cUEsH
e0qvxDKDTwhHuLKu0wgI4FbZzRaynl4F3+XhH5VGru4soY+i2hrTslsU5qfWq6NWJ4/cgSTzk/X7
GfU+9HokAYL/TX9qjcSl+m8VgaitSemUnCZFcO+DdtjZg1Zu22Sd/vO9FHVt4GNyiVsUJdW11rM0
g9+EHZN/suki4Lrs0N8ZHgR2TCXKX2/MLGnSM/KiKj32nCucIWpaMINU67Mn2inOm+07OfHTtjUx
dJXiNjdSrNkzwNTez77XbxTP4/MvgBtgOTq6+Q0XAPmR5TLIwEnfaP/hUiKHP7RrP2uAF27r4Qbc
mlgLHr8Ajb42t7/c0raRIJJfJLbFX/QXH1SSo1yqdYwdQAqdpvPr/j46OkdEW3G1o5FcvUDLJmt2
5WGo0huvhRcrhjh7SMfCjj9R0MIG43DSOIRmsGZdvZE8iVTrlLyIJCvjr5t9DTXj7iQTH8u9p/Rt
j/OR5SkZIqg2dLHjPa3NYhAOJEVUvS4Iiup7nGxrLAULUYXHwS3IO4yOyFbgKUDig+Nk8opa3bkt
5QLNF27RVxF1bFak3hYbWkhGibtTPNqHIAlp24kc5M1v7hVRr7LrSs9Ro1pMd5haDEmXwTg0yd3b
QIpU8l8ZHwbUnZYEe0uZ3L/8Rsv2RvJvqw7W0ahRvYfQYUyP2miPqHY5WCoJ/S71Sq+WEaUK0pgy
aVFspzOG3yo+2Re23nucPzZ+sVnPWKNJlDIsoat3spgWmCpVMuUj08stiIGrk7ix1ZyZJPDNb8jk
aMfouam4UceUtBtPwLO5+jqZaABV/soGKIBC69NfhaedN2ccq17BJdh5rIWCTNn0mhSeDwJiR4PK
1fCoK7nAfsxHBNnZ1OhXbxIt061U455QM1UVGRLm/KAKZuWE6XnwlNrRAUwHoDVQp97VFBQ5fGy4
MWohraPTP2ZkzG1sbpaeNI7jHFoAXyXAoHncBp5/iUjKJczWH0U2tzOnmLFC82diFqoCzbiLnqOB
0N2Sl1xJQwHLhc5O/gK1GARtQXXGNmX3R9OLaCUnDX209KmSgZgvQsflC0zHM4G4dS2LjSNdpA5J
o4zWj5qJecK0Xq8YTz2sNEcCElVw3bTHIj/EV13Pcv5TS6a1TiFTw4lP4jvH5oUWvdo1XNkyT2Kf
FkSniGc5PtKM0m2j0q69qWkf6Dun463Ms4Rddco7lAJuxSY/Q5+POXXSrnK9HST7QULfojMgBNyU
FEVe9fXU+XxS3tI/971IkgSqxUJS96gu8Rv2v27e8iuPTo5QLnaj3kFH12hdvfgmxodbK9277ZdR
W6TqXx1ef1/zZMEkPLtCuIjHsrzAKvlhefPUKgWjVzuaNkpwPaY8mr0LEkvBGJGy4vA45nSEqOiY
Rie4fcKZ1+yUwoGBrHrs3r2G9N1rs/MorVBYtWCxYVTKnbVZvnTXMWWR6HWlYk8/fgv5cmizqeb1
r3IzQQK5U96ZQeZ54zDQqKe25gl/DlH2Q88hfj8M6fqyLs1XJQuuBoigVFMHveD63nafDafkehFt
asoCRmvNZ5KXraiK104ioJbKK42/fqEHDoMExylUWhMwRUasiQgwwTipHBSQXpNM8MDthWMSr3yy
v+Vd4GmqjxiOjdCPacZfNpmoH7UgC9WWsSEzjc6o3Cka69rvUn2d2tYN5KwZin4IwbxTE13KkWdd
qMAkbp5y8WJz9gnDLfDbXB68WB8+3YBvgNlRUurSJcCjo2ZtbcMWVmMJx+CtsnpgVLCVtsGlCcrp
mi7LcvmwcL0fBsd92GolyOQahUzgS0fybhlVnLjNyYSarPZIYoSq+t0vAu1e/1ada3atiPpL+8++
FD85T1s49+gvfgNH9iRMuTi8WZtdgbLg2Uh1cNkqHIqYBsepTbFpjCkTset3+UQDriF8utQSp2XH
+ygPh6zroQBixvZLRMuwhyRgqDD5p/t8pyLp/xvuaz4na5SzW/C3uwacILu6uAJwZ1BoSsQjesF7
XfIfFCtUL5EGjH1XUvxwgglnPDIK7805qE2KIPBVWDHm1Lf4A0eRY3p5quTyA8PWzI8ejAHr9Jcm
g6LWSEYXfYXI02jEAri0Zk+HSra2RcIL2vMa5LL6458kNN+kZVGm3t1zKW5skThZQtVLwoQbww8S
x2rvDoKf8a2L2+fZZ7fsaR7OQoLO25ZoJyTdfIC/D8Tmg+osYBSBa/DCdrpxE/E6Fow3qvb0Bq5P
sRh5KX5yONEveujUNAIhpt0O5lmC8TEoKqBT2xPJoEJWFHVSYDTeHJAHLtCLkhZWRZXLrws9HgtO
YsJOy/9yJZOhLR4GbgyIzLhRB7jqFtuOIEsqgxRLrodObWtRcgIpLN+y/lS7w/1zUU/EqMs8jUXy
H9/71SRqRxPvNypkdZky5v1qb96e06Ut8uuUE+wOZdF4D8J7J1cp6XMstVjyuUK3DEmlxEeFdEmh
9HhHG7EF5voPXup9U9TZz4txAKpLc2Ot7yq5LII/Obk4rWxr/Q19d+4kb97cEhagP2By+2KidNKx
+aApYh9BAdYtohETb+TsrMwc4A/gLYV8fyJO5m3Cv1MrxRVRtwDe9I/QPtXzE3OaOnIWzhTun/Ic
BYHYPVaEjyXLoIN0yj8AkwQ9J+n6EasR5VUJCdHpOs3/Pb7hkZ2yFvfJTI0MTyu+svi29offrgDE
4XSeWRh81qaU8dp6ER3lDuPx8POLS0vPxi955ftVlFp6uxLAw/kexp/W8GVbYicNYGPeYXHmgGHB
eyxyqeINQrRysRNdkXlatj9blJVjUFCvCHVn9CVNVW59Bf+qK+UlYdpHcrhDsfXhqORd0qnOpEI2
7vP9whrJ+hAkW11fIL4hLwfWTfp2XHSfOurFHWv81xgLd2VBKZLaEcDJ1yEu7tfpRDGp+Kadr3Hb
id0L1Hvgju7mMOPh8JerqehyS3fbnet1ZpRU54ORQNJgadKZ38td42RUKBdOv0L47ax4UHmLoSOb
dmdq12vZpJErcCFtUTJ6/zL9O+mJhjdmfiS3x57qLY+SQVFcx4LfmCwOfz4IZYmAC3PIGtPLNzXZ
P5SYOFd0QH4LZBoONcjXdLN4NfYV0QOjZE666rQhAx2/MGWTph7CYabGNVlCPvDMHDMoZ3eqkmj1
nh22gM/EXX8+51aMCRiKVj65WeH4XiWF5NEB3/YootGGAvzdi4pDab68bNR+36v8mChc6vKVyGhS
B6c0BdnhEOJYVI9iiwclnCEp0YA+h9xFfh6clcHGdbbV5RNpOjlcZka4mO4Dn7R+fbWbz+lpjC8h
M4irlX1TP6w3mzwiOc6adtDgfUnwS7UXU24qiza/9sfEEYsqcq4iBJu9c4qHHdhs3fY3Iipx0F4r
cBqoZHjRTTPvDNJIeIXYish4qKnNHADL5DP6D02rN5+3k3B/TG/FwdsnwM711jFny71CqKQ3a37I
UPmVyKTBjZg7CR2Yo584IkYYWFYUHGCttiv+mQvpt3CgrFBGHynw4vucdWawvtI2KC6wbG29uq7g
BcLyHh7flhpdFjQoPshuiZMUIivOhellUEYzVV2tuqxnFzEgXmndGLL5drmEjzEVegLr9hAzaSac
ZzBCu2uOzPB8ermnbQFutRj1FU2e2VXmb5fXFxteg8RLYMIJcMHqLRe4JhSIRIJh1RZXzMPpVfxr
A+yMSFrhky22JYKdk/n5Om3clQrg/lLTDUqhA2nopGe35o1+kW42f4zk/MjbY0K2jzPW33qaFxDN
YMyck6U1WvkzIYoWcbQNOrlHhzo10MBBddBNlQDp6Sru8t2CwWxl5dASzog5kBX8OQR5J+NMI5ED
GeSJ9LIHg6mrGENwAbEP0kUBQdMU0MIMWj1ugAmR0p5aXrlNugodyy8qMeEGtAZs8TyTZ9j0eo52
r64RdL9+oOuz9Uezd+JxPfDw454iwGXqjo5bJ95rNPLAqA3oHocdtMkKCjp9dkCVRiMXkUjU98iO
//0+3dDKfXJj43sJnt/N9mDem83EtoBiVde4i7yeK5NMhdUPvKdKEefVCBRKJiaiW5nBrSmWNB6d
uWExn0dG5pWjZLy8ZkkZpU4jo4i4PWXAKLk4VhmR+54vMY1YviP03/W+Co0+i/LG1j5UXq36Tled
biQ+IoerZLzbsjf7qVb4Rqvy411/gw144qsffflutVnY+iDTBqz3pSoThCMEWq6Dlpae8smx7nkw
fPK/SJYjKv07WZfgZ6Zpu7VubHsm/raDeyPmsYvnZKI2gkso/LY5gS4razCtmGhWFMpMYTGi+pVa
DloiaDtEwrAYq8zpl+vXsZbGJP5IwxsqQyGk4z0DfCT2hoNPO5pKpbv4miAlmpLmzQT9TLi5E6q8
pU5dSOIE6Rnys8284K1KSEiNvCQYtd22+8Qi6t5d+o0fCgVCqpxS2L+yh/GXfIVn8KcMGtWUqAQk
Jn87LcrLQCVqKDA8fQYQeEOgoeXwwaes3xnHm3JJ6XW4I+mhHWp29rXPDl3cTgB7DqgK9VwPxiZd
P8DsACqiiIqucMQPCp+Vp/gmKCQhHURKaMhjRT0Sxzi0r2t3Yj/CAh0njZ1KQLagyqQLxbXAIyAN
7PDZ5J8GokUgzcvqJ3lLfMR0DwVlDoWVDsV4M5+ImGlXbbNbwvc92DEtERS9xu9/LTIpxE8TKSbo
k67YirRGZToGQBED/4nFlsmErO2ahQPgHufw5DurUgT0Cn52oSy1s9msFLzsDKQiu3aX4c2xJyQF
r2doJNbqgAJxsSC5NGfCyR5o5Wy/pRaO9uHZrfIEguWkDvsH/5Gwb7KGcviqYCKQ6te1dq319swc
fZksu1mx5K4v6ks/sbFHB0XtaQUOIrmQHqSyFe5PTNxHB4ajFxxotD7l9iGx4JxD6O0Dv4NbWDZv
9PZOfypdtpf9wFCWDU50vO5YmXurp8ixM9BUxPc51EZgAgCSoTVRjfh7PRC0ejAyWDLqg/z5FKj6
CfvFYyp3paOp0evEj/ieNNmZ3QPZck4OLnuUfwTj4BKTrQPkF/D4Vja4GJXxQ9kUma5w0c2r1gfR
Nh1l2aaE5nY398hORFaZohX74Y8pc42tq6tckzoftuZY6hJq3VxH9MERXERKCjxSVRs99VLBQXqB
qwHYROxfT9mpvq80wzWgXuT4ymtOvtqtPAwmCQ0VvA4GaVYi4IHAHs/oIOM1448AAXuGW7zRncAe
2AMc9Kqgq7xti98y1IZynvly1Gj02QMNEnfwo1LJfOpX01avEAQPVmFlUXZxK7TpxFahmgF8/yHH
UWaEKuCZj3u3k55hd+GeHFIUQP9epdp3oUEuF6tNZVoXF5ZUBXyCGzY4RUh1hDvHlvnJxeC48KG9
s2AOh6V3KoffvlqpVl7x145x6YYN+OMZqjqGhFsodquVJ5gjohghzNSRBf/9oowoKk9UotmZnucw
L/13RisF3mv5Ozebi4R8J7bHiJRYP8/4OxQIDfXl2XbNxKgdFN1H+suCLQ3rRI62e5du3yDhSq3S
uJHTlGgKHR2w/bqMpdExFISXxGLfndCnDZ99IoEF5aicv2WMNiPxtcx/flgCIh2ncDKGtDDITWR9
XxCD8/ROU1KtQBazfJnz9toinBXT/+qQRZI9eK5BM9vxpZSxqR6ld4ocZ4NW5e2LdsPib53s5PlT
F9WcdNp+IWMcf/nVZD/gXl9N4Lc/7PTg14kDyMPdB0NhgPYNw2bBpI0n5liKASFR/4G8Z/kUkrum
d4HG0CxxPRQujVPbwv+Lt1Q8hk6vxpx/X23uQ3T/KFdscMekD5aSb3FLTHjcJA5WN1oAhh8NnWDE
MfBnHqnfQYWWcNiglbuBHv+hV9HwCwpWQ+WuIoV9ZYWDneMKm6bL7zjYbPU0SmgowyPx3tT6ckKH
/i0wml6XpwuVehnToz09G4PgZFxSUOuDe5EptMhKUWB7UMOLNptw++gUsHBDQdVAhcPCNyGUVkEi
l3c5OKKFXgwjJ367xfZZB4PhOSqlNzjKsZ5MEOJmpxlMjdNs+xYs8j0yeZ78A9pJsH/IjC4P8YRb
aYMsMjTn2g8Qsi21BIFFrX47+6elT36S+tBpfTVgAum8e6MBqSgxVQyuFK050aN1U5v49Ji9cmPJ
9lmKcXcdo9sonwHfnkjePyEvLIMK1g0BUeYOZH6dggEd7IDCaqHDt2dDh6W7fll+oB/uZ2MYza3M
2TBVVJCh1gSPoFI0gULfFzLAZGeEgwqDNF+rLYoQ3oNzXROqNR1cyCeb51bTk39nITh+hPXyWPT3
M3aPJZM7ScLPuDPh84mKKsmz0j7aKWkY931t/bZXOkgPaMD3DWH8XF5ECLlko0ZdWI2HJHwXGc0Q
A4Fbck62QaLWwrp2vzipGIQkvZ4J7qxXX83wNml/O7IXnlr4tfBxKq97GNe/RGmOZYM/DP+M4XbU
amefiCSXewwKKGkAB+9KT8Yw0ei0QDO2yzvEW5IugoWSIRujEJli2vvndSMs8dt2gIKffrKJrGnU
KFGr5Ymv9t1JNGoouxL6/dZl+TYf5+9ZbcN95qyL+C22KpgPV/+SImIXVjaGT8jxE6BUtcJH4xdy
YaPjgIlTYiO3W7R+sgI74nPdzsO9/mfUpDdZP2xIAuyaZFlQX8AjAIHHtvVqTwCTxPQbd9jtyfvP
3z0HFjV10Q0Ifs8CazvZSsFoUtSx92u38y6FfV5YpF0BMP9hqeLw6LRllcDvmrE0budpk050jtQP
LZnLNggREeiSQcF08HxlZP91pa75JAGQsJeEX23ukbukQKej/KB3joKlUr+v5jQPI+oVqjk8lsEk
uqre5nMExE3bEJDWoqJqB71BaofLAMRKKxMBvtD1r3c04iZFCpD21JfPxAMHUQWh7mTy7jkTInd3
DdeHiQydHW/o+yoY1H3GNo/qDrH7LtaiTo6xQoO51nGKWTQjxbZdEkNHHHbJucGKB8FbJrwn/t3U
W2nlawH6HCGy5k7nGiz5DXZY5soPHZqeBuVmgsoNbJR6uDB1pTCm4+2XeVIZTh4hNpbm5RiDasFo
NQn8sIOzFP8nsW7yoWzBcqQjs+gmL7DHO0AJ1Hn4NPYENUuCoQIj3huNxn4QapHrHLwEHFUIwsbn
rQ26CfuROGIq6A1stmKTFufdQEyI7ajXLv6u2PSYuCU1v47KfhtGPBb+ARwdlCMr0hBt8TPmOJbS
17ILmAdCAex641g9rEvnaYNsqwajCXLFEKATfwlHW9DfJINZgBz2IlStAe+rt8hA1ZksUqzm7kod
kY9H7GbfGsxEzUXQXk6Q/bDRif5cJEUjrfAQl4I2iYOkOcT3hV48SX571gX9ZaA982eXT8SqsXH2
8NROVGXYcsorP4u65iaBzdBybcRxEa/xCENGzslouK+GSe29hNoWw2ji8JkU/zhZx4Kh7lC6nOiv
/TugzT2epPDyHBuzQFiCiAzWg3VA4x2NFk4kqmspx2eAHfz477McVgCxKbzsMdgIEBEVjyX8wKXf
31eJObH2nFAwcpOyGmGiXxBsG8m0l9Q/tmj7eh2Ed6aRsuxsn7InbXKb2ur6yGUyuS7cTf1PiTAP
hnN+YhFwvuf5vgM7MM2EPpNZDt33dzVKUSSxcw9TTM9f/uRPCx8RRr96IgazdAdbgbPMtzO+IW66
cnGUee6Ki/b959lTS27mChY7Ez1ck73wA8adB1eIoTucLihEiQ7BxvJX+b/yWQHarjNcFCeZMDw6
y0lopk5SFsHCVV52rSEg1ngkmOIB+wXr+0LanPDF1f2PBrHanpjTUM2wW6NPk+yEvy/5zv46kkEI
n4AeT61ENtAVcxueWIU3KFZx+V3BS0961Q+soz31lhbi/1GdtW3w/zafph39cfjRBEmnDnu9R6Ym
ZN0vtvKyBz3PCMfRNA3EVNEgKVlhgYwYKWzJiREk0lK7GMTAfz1RDAk9wgTq6KF3IrWHcGTURnAu
ijrWr0B1K4fwdYHk7MuWG0l+TJ4yzJVEVoziqL20bqCZvQokEg2Jxng6M4tmsi1ZeZ0sA81cj7rX
ZZYwq+DS3rA7ujXlRuUgVXVBhoFL835vUeITe2jzG9Xkj/162XTrY3z3juf0bOXv5d3/8YMVQBXL
HZNOoXnyzBctocpNdoFlLoqI0f8Q37Vw1M3C0mX+5MHRC0BMZYRLLdGyPgUw1GaPSd8r//cEvsfZ
PLPPStvOPBYXx0xcnWaf+Xc+844OCxAxXZPe/c6QjQtkyazYH2G/VsDRO8VZ4YmMHQ5tSGV2KowQ
/cbkJIljwV+XgtSKiUA2X954oojFmWVCPlfhqSX0EsBB/h0Gz7e/LbWJEYOnHVhBsiw+vE75g04t
2HbvhYnYcMwoGYxocP90haqkjwxhqVNce59KM95PPWW9HFkdPEABi10A3HQeBt2XbK8WDazANcz/
Fdd221FhBABkfz3DmBNSetn845J5MHy1IIBN4ReRV1MyEYFmN8VnWIU+gduOsvDI2mhf1W4dfunv
cjfjS81gCAXaBHMLfRvvAimVDL2wuUYuC8cFNBN+oYEpxhGgP0UxPBx1ZvYGsrT5bgZsA81kpgk0
m/sjRT2HXDMrGoHdFYXCShUBg3YLgOUe/hCdzUJ8pWxqxJYhtjvprvzb9gbeCDjachpKvaELDYE5
woXO60DYK4pywQ9fI2FJu6E08ikjzkRwMlTHfKN7Ji9Q3XujS5B9xOj6cHP2mpk3yoAtwBCnK01u
U+JugjEoWMbLz2vtfbeQu5IhRd2QCpPpme+So6d8CK9GnNaGTokTmbXorL/cXuXp5nUSl856o20U
K+fi3OO+CWA8Cf8BjxrwkXQqvhFyQW8ZyxlEwNR8wF9ZfruEvAHwkxp8A3cS7Z/XVYKoZ1n+WfqF
4NxVMS75VZjjyOWr5BhakAydRYRQB6rC1JLDkT8SWbEBywhYpfABE1FCSeGj4/gS2mqOKN07NZDX
WxdqdK2+ZJr5GtPxwNh3dr8JxoXTX3HPyi+NULN/uZKXfl1/1iEks8V5oLrgaU6yghbkUdg+boet
NAqXQTrmH41jQW57FbZlJAzC3e5j0wiVSHwNg9kGSFSmNteOF7Do8YQNeUvc2qBb8wyiZOcO7mXS
N4BD83Qn8OdQq3GiKlbUhs2o8O7/mGWLE/kSTtXl0fN7eytwaTGNzyfjpam/ToEMMMrToAc17kmB
qfprPU6WghIMrcr4a+0SfrBQbxdahYryZr90qLMqsGFdJYk5nZJNtMklYzNNJC600vdzVgJCV5IO
+PYQH/CUdQwMjd39Hjbxo9122FnQnsVltxVHV0LMY05xZUpzflGUgrZ8ps9fnTyFfmBQoG9pKtz+
bmbarxxEvr9o382WqbzWTHxCH2xj3pj+Q+TPjHd95IWTgYjDmKMvJIP+3Ne1RcCO0mj5lpouSYaE
gh9RDZDcmxFo932ChAYqM5ulJH1L/w1fg1FWaZ13dAS/1SaaWvzAYsohgLtHzlZ0ITr/DoR1uS5Z
5GJb91TO/La5WFrxE8zZTtbBSb15n860MslF87b9/Kt1OBQZvOL+Nj3OQLa7gHUmQ6cdB1BscE9k
/58D5gWxMMHT9WZxSQZUByWvB8kWcO4+r5IB7ueGPhoD6vGER2w7+4OcHDLbcki/fC+L8T/ATaND
92CchHSkpcAK7AUTIGFweM7FiX12mDq1CipM5j19gKfAY5tjtO9KwkKBL4SkJxm8CL9P2/0amx3w
mJ7uUOw+PpWT0jZGm8JL/r1oNVriNvUXwZ1ckOnHrsLiYDv8tKdnLZ+uSwjaV1h+4Awljk6xepqr
GKiLkZ206quvZIN5TwMJ3mg1uy5rxHZccd3KrOxH3aHCMX4OnszyLkA6L01PdImMaKXxaGqduABJ
vMIjVR4StEx+ea6Fg/pahUpFno10fxTLm+72Lx04DsU3yxvlAXl/GJzaKMwXgBX1taiu2mpsB9yp
Hp30kyMOSlqULja3vpLeYDJNC46GPrh0i4N6UkUoYxzZ3MGtDs/8vk3Ff+KDAXIjHgIKJwmywDyU
PtTuxnCT51AO4u7Zi6wsEK4pxLXoJ9OHJLKPci+0RNGQAXa/x186cQWYt9wewOpA2OX4R4cvBBTA
bdXCjvoJoOr7/+VviwCURSBHURDYpnfKJCbvjQ+TpEj4dGjEBhGqG+y6fURch/e6dV24oLjgD2al
xhGzzZCbPdL9/bXniBXulzClSKCTuX81olU6dJhV99dJevGcQMlDZ2s0hiFTDKC9FtZLVSaPxzYv
sXMZMMlr7mcJXSgZsMlrqtcu1Vjq8Cu3fgpyhsZ+2Bt49py1wnY0Ou7NqjfmL7muVVYJMWREh1B1
ndZIkRUcIkQ+wXmgatH02UORq8rET+d58ggGF4u4EfI6D2RggpKLsx/lRBSl4yM0XT4lYsnko7hC
etEOg0/7yKzYG3UYhBkB3u3YOKtsBDnExecMkql+beFOAzFf87p0Np9leRgc36L2at9GHnZOGIm6
NWGESxgGMP0OiYLJECbq+LdOvZBPX6ujEJsHSV8R9ZfU5QCkBqF469hFE8ZHHytEKr3BvTtPBL94
fM2zcZ0Z0pZu+T6LAesySNE3CyfUv7vuJkXsCrkJjLfmIEZ7cUoFaCtTAch1C80/IogNZZ0Wr8t+
J4Ay1NjOTYxt3qst6xUw+A0ViSF6KWP+8VpHXKJFYk257pFcbVRICZBhdQlGlTQCW/BL17x152JZ
UCGcV49/dwqKrZDM2dJaYGGy9KMee1VL3/bQM6CCJLS7uD15JThtLHYezmJC3tk8FQdRDM+Nk/h+
w3ZI9xR3lsE6HOPCZ4LiC6Q3C3m6sl+e5eF/lzlMrm2d6s89QRUtQGkUQgRB0Zw7XPmJ9fM58aTA
TV5CRrluT3lVcBfngQy4hDslh0cdzQd2ysiOSvJSjq2sI6JorGMjMdjX1aOPlZ5V20uQmHo2j1N+
bOJC1tbQ8O0xq+JfA+V7yIr3wxUCrIej0t7GkcIPx5wyVKrbO87yXyAyW3KnA5a7JWGhUHx9m9E7
Am93FN7Modpi7QfOaTFP2baFfKsznxokjB9pCBYnqn983PyTqhDuukjF/8YCVHCH2isBr52k83Nf
ApBdZKsPlrix+R2/SkCBx2LdzN0vxpkphvad2y6+uFuNMv9JIsnDgE0tA8V6VEqR75wDE5a4tNpC
GIY5jeQPvln9YUIpibk1TV4menj4L5eq5QICBsw66LtxxHqakB9dSHEEW3QqUimz79YVzT5QaSEC
4FwNQ2Z53sGtQKBPa7ENHGsGfu+KTYGK8H2pG+XCcHEJ8ubc4wtKWmikjrpPVksplA8/aZuAFfTo
TIniJUKhM5sBBWJhXtMhVcqNsfUoiLiNg2L0jMVkjo24zJqDiNzAwMAUouVWbjv2Aef3V8Z6Z1if
Z9MUj1kWD61b89k1L12Q7ZNrrG8JdfXOpe0d3u1jziMFTImgSeYhzGP3233HMqDBNWAXsxGiPLuA
sJa2Prrey3ENSSmLPH7urKsBJHK6C3Hlb03U3eafJO44fSa5fuBNte1X/sEk4BUwmCsmpe6gIl25
Wd3FdamuwlyYVPgwZul3kHkGBFCAVXheZu2JlsYBEvyvG7S6VqJia9L1y+dVleZec5WdEl4c8vqc
EAm8TEzjBW7UXlz4QY1/TsC8opua6iNzezZe7UJoATha0fF3DATwght7+m9iR+tjmpoLZledXZIJ
Q+wgVA1WJoo21OCpYRXp3kBpKAGMI/oWcGxFZyzRHQMnJXqcK6OS5LWLOrbh40F6uxpQAqBXlfY1
h2heoIllUZLzLOUlg1WIGyawjYBnPfi9spcOqufGIQ8D46Cr6cGdmKD5ogGddLkeWjJ4RRsCvdev
T61PPNXoMuWyVjB7oRqCxsXmeKjvMjZIWD39G44p8MSaFF6ADIKi8V69MI2eWC8MDdwU/Nnequ6M
QIwFwaiICJuEUcxpuYXpY4Apx3Lo1jFQu0tBISTM5ttZ4qab/GiUEkzYrJDGanehhwAvjBgEOuq4
jrEfWXsFGjuRCH51h2n4xLC0Mzg/ta8Mi2JqUvubFaUdJAXd0NRDdqJ1XdwMj6EgijyCYkVBm3DD
B9od1sbg41GK2Qgz+wy4OWJPYerijkfgnysWOm5JyRVEu7e6BxI41E3XhXo99LMkrJE7jxYkCxhC
oJ8FPX2GPVrdpquaTvHbKRIhHNfDx8Wf0T3N06Q7JBC2paz5tJYbVwKtg0eAfdaKSFqPZHSlR5i0
mpS5VNxgQBQxtsFzNbaOKu/+A6DPfEqRln8N7no7lYoGbuHgy4U5u4bODHPMscu3LHnndtec5ow5
xaq2FMKhG8kpfKclCfU/eJDf/U40QvraMmbieuRhtYn7+L/08SLy8XYObwnRTEv2X42+1cL9djTn
0NSfG8FgAgSNFjEiXpJcTN+03nsKKSo1lMiA9EFf8PdMfcfmVCSakVNrLWg0DQ7Q3HtTbVnTxYpk
CHbC66HglHB9keIQqL9tMaqySeAd47aQ+6QKbEY/IYVW1IZbXE7QNrsR+La2khNx2HihXB+uFW2G
ZlxmXWTrn7lXGRwyYE316sFDZ+PR124sz0l4+0EQQTu98pY/BFuHdxQuvd5+y4BR1jv67hSF7Kod
/sHdDyANqK0JJ3hoWrSrKF9rhA00qxER1ElJ2KwDc5r63loJ30BaQrsIho+pER6fiaAyN+28laS4
Y6JV2LCu0Kbk1sZhzc5N5WCd9Lhbb9pd8sRENSuj+7ZG1Jax3a46GZ4pkjA9YnmPLlYwLROQs24Q
LuHJ2XYiOLGmA36rc5zeqnz+Rf263YsewB+0rLxC2h1Ot21FdXwpWd2eT4gp2xDR1JLlCkcjqera
+t18ypCtItWq5Og2RK7ASRToqS5B5uBN9Qy+RuZPZTgvHGjIfL4V7+dGK7tyrHfuG/odyWyMN6mI
BkWPMG/GkId4uySwznajKp4eq0J27hHrn0B2MsMtRJ5NyZopdMYAOevK0/4mnusft7V/o5vErVTz
LAftQQWiOR34Ws2wZHtxXKv78bK7EZXrgx3XGOwKV2B05QAhf25EmZQ0BKtwzeEfLAalkjSGUQs6
mNu5L3YUWhTt+5rR9dATpQVlt7oUP8DZGVB0x2CPzHSNQPwiRVwvWPswMRACn8WDdmM0iuYmJGyT
ALLJhnPb0171guStyjNYn4EXnA7DKD+rA778dJX5X1GUNr1LJJg7oLY2dj+BDz0Yd3lkvmC9uLNz
zMrWRN5/0lTmxiXYNzIZDGFsjjVeE231HDY1H/0tQa/NofXruuiBaMCSy7ifotd3pD8RXJ4gOGnE
67tJ6hIcPBUdyRbEE/OZKqfaoHQjqC4x+E4/iBX7KKhhgdV/23/93eqYcQF55DGAoItz4IAjnyk0
zRojoBufO+FX9aT4dELC4s2jfa3larKiMnXwiwlFdCchfLlWkzXl+QzBF/1Qt/vJG43ydPZahIW0
06ME9NCzzUwVnIjWi42or4ht2udExkbjVStl918iUy6psieWw/JRcTiyGqqs9jfFlHDA+yiJL5Pr
kYGFFsbbQVM7XBnz0i7FSIoSYAfoYI9GXPnJeD1uCjQGe6jbrQMUyPsGaXncAFRLFMquM57IVh6O
kf8VRL87fWLQd+w3giSAI3NfWFBPV263ntW6aukH+9teQxohK+ZJCykmbllWxFFIP5gm6O4Q6hUk
99McRTKUeMLnbnOZ/L6nQAUSKHAfn1csMCKnBaCHDGH0tv+PdLvWkgLNTbM7tHtmPs/3P8crwSxt
09wPkOM+36mp7CjnaQpLq176UD6mZwZRPk3lRCgPI1Ih7GE/tVHivmqflDzrYovy8LUnKpIdK3Kx
33jFgdt9PIrT36k/E0Wq5BAYeMlwEKqRwX0ewSiF7OIDPiWZEIN+/adCBQA+PJRh9MrfeyK+h0yi
m6JqRDySYPUweBpEhgNhSXs6AC3DlmDY0eaYi/Fd2LVlENE/xrQHR+s8FIXg713N2BqR8lftM6mj
x17NNHwDt/pmUnMp9k2ucZXH+L5ZtycrqJeizqDLR75UEeWwiBCakIM7+o7EgeI9N9Z9TlqGE1i0
qd1HezwHvHlNJUXlgUGkvR2nowbst9JbYCDbnpXng+SAqvydM2aNcfXn4LFeGwpzpURfrTsR51oI
QIYL122/NaHUE0p3yAEHE7MsKErnhRLn9RHGjPpfL/HUGT8DdEKXmCr2duG9+ZG8zAs5agjjXqOh
rWSkRY4eEIZV1n5mXX2xuLcTOWr1loMAv3LN4ZODEUEG01/n8qLr7RrEWL4KA1XkREaAVbPnZ6Uz
Xj5uAaOluddn1yCHqaH3WP6bQ4lH+43+JRkS9ndPodIdyv3MNHefmcKQI3O5vnvxXBugDIoGPoOy
JrcKPVJpfQSf0kGjLpAkhIyjUrgGa5TQDx73vKztFaqBvCgljiz+6A9XgSj6e4tS8cAV8ZAQ47l9
y07DyawV9RmMAKMrpYrP4o5Ggb5vK98UuY2MnCZ0CP5JVb6Eycclysg0TiIIMV7C0cXfa0lM930k
rAHcJ/aAZDl1H+Y/IPSMnTNQ3IEcKvEC6kgp2jpiodiehzznE36DideiUb2roHolMa9gPPPeLRja
oLonLYjyKEhGkwms5TH1O8PDUBlJEp9pTa6Co4r90qwCMwHg5yOufoNHb4X2W6U2d5z1pcFhFEUH
J3CuDUG9wjPsm3J/8hXi2bu8ZwUVEd5uPy90lK1xXNythJhu48C3Iw4RsmF4VC08Mp6xCb6MIvSX
Z11J/QGlEt4bsTzHQl58/MWhbWnqVBdGQxNVuo7l7crG+UVRGwvCNoPFdAxzcpyi7ZxdYGBff9Jn
RosTDt6ksOuXZI+3RDFcmyx8h2pzrCgSnR4yw7BK4SdUY8AJp3DHqxTZOplSeV7CSMnxMEOIlYLf
bxgrilKhr44OnUPHCUlvvL3KJQ/zu/za4e0zc1l5cUgAs8JP0Fv9C88DU/Ubx6xsyXnne/qedRNh
GdmIVxRMg3Ny8qXKVB3BIt7WwKoMfPpg2FQ7a3bunYYRPWGUdPNT5FcRLFl5D0xxfvJFCvbx7h23
MggjrS63DeRnFUOky4fa2BXgwDlTZR+Va4aqSHUumgMEh0iUvr2u+Qz/YNT3ntVhfrW5VQzOInyN
CgGNQ7jB2lfjL3uiNTXmRz1q5D1j4eL+7dnSdCSUp9WB8SqfEH6nmy06F/XK4R2KslXa3f27a6Bc
mNfoOJS4Z4OooWr7En/zzubJxG6OwI2ljfTPvChH8dhZKP218xKJn8HI7No9HfvQG0ZikO7sVOYh
uOlbikGeG3q/ch7pdsSMYDz3L4IbsikJoLs8Y0GKb7t/1jIA9eb4fA66xWSJTRGtLhugSQ93Eox6
w2QWKWdvfGZVbvcrFmFHdxXvCKiutfHLsj3veRYRmSV07iZg1lMLe96lXrqFCavKFomF18MVJDVW
C/OjHYBxSRN0SWKNXV7YTTtLcA+eUfJTh89VFsrm74NZdZKUMux7rMdXwdMp43rpt62+RsiOA3nl
YHH1i+QDqbA1er0AOkvC7NruEk/oz9cK9hENkgWrFo0Y9xyrL+zYSlmJwB34AjV6Ls7YVue0nYCn
H+mHUEgKfPFmB/+wSyr7Gp3Tev+8BRL32JgxjBxEAJPbpSGK+2aGvO7g9mTsDrDTcPzNGRdmeFJ/
qj7thfivnMAkMQUwoN9k3UiW6uRTrbAep6PYW0CsZUaVvnNNEjTKzBbNXhoAm/Cbe9lLGCvidnKW
W9ieMWp7LeG+frG27DI7d0pYzRp0rJUzUAqfNlLTHaLAagU7Vru225kMX7NOolcS1niTQxaWWpGn
igrI3pqaGyJvfXtJm+REajo2BmL8igVODkEB/pAYm8YKMPEYxIUSBJD9ntG1IV/bTZb4/KwujCAL
QNRxyVLKskPUHfjziC9iAmBUWV9P1kbKZLNnDMo7UCzq2tDz9WPNZdHIR2NSxMBeX4BPcjSPSCz1
i4zy/7FEpMB77B4qfOuffSk1eePPp3o7kMu4BlWzdXJN5y9mAyyk/5+Czgr1mVytpddsBq5B9XlF
xby5rgXxJD0TKwsO9b3s7FCzFuZVppvak1vR6qIJ991jMvHRVn8aJaIBwL80pT3m4lb6Fq73DwFG
QN1iTMqHRioXtj7Rk7N7jj4UMgj13yO8vNNw0tDsWOhlARfZa3Cn3Oj6QozjM5HUSfbjgQbTcE5q
mTQR5N1CGIFHPbWNGu61ZnngXTJRwblT8FHLKmJmSllAOGYDHpUnzPSIuFzC6P7CT2cDubU2CPcN
mwcTW0SOSxCN/2oxoeXF2kq/zcktK49KOQsG6BjIMNX5M08jViuRutLNL33oUHQibeC5NXnUcpep
6srV1my+dC/t+5IaKtbAz/FGQT+bQXE1pdJ4SVwckceFSjQ0yi9+EDFtweat+p8Qp4Fcy+Skwe+9
fSvbTfDjzScFwivq/Y7SwaqAnabQf9EMgAr99CqSBY8ll/Lse5iJvwqix5VHxXtAGMqXAQ+9LEuH
qAmlBofUbpxs6+V4M+InJpKqyK65fRdMGT2KbMiPAocNoRnfFa7uDZwQI+90b6ljqOmX7iIBWV6H
Mj1RWfwMj01L+kjhMObq8U42zjY0c1YOILYyeldewXUTcQyWhcB5Q2DIKClk23nm05IVAb8FskP/
/mNItQt9HpRCECtz266hohU23/iH7IHV/N8/y8F5SuikG6kBNJskbrlVRSJj8gDH11r/WF5KYzQS
ys+ZklxHAhsBfGDLFcgub2W4WXCRE9ozrL4bXBesg7fa1Yr6pcwNMOHTRaIPALucTGPzAAxR/Kpy
CwhButuNmav7VSj1NVc6Uw1ptL4e3u8KlQ/akSs+ePvlfLihKO0ci1LPENGGN5QW9xtLJDtY4jqR
1XEa2A4gJgal7bK2dOdGScqo6wOqkoXPJ5v3Gu/VBwjMhRGDpCQZlh4htzY96Ky4sp1QmvVInN+B
42qMONiWGR3KZFxXyms90ZNgGDM3De7moONVfGOAeroQvCgmK1nsy1BZLpbd7nieCJC1yAX7eIkm
gBtzN3U8CKUSeOyqQUMnq5MO2NSHnTF0DhiYUdZKE2XI4m+LpFkHdPvFCls+qKoX56tRt3ZcUaSQ
eeL12tdBDyn4bPUprrkYpk0YPMja8DlVeIWiODqu224lm/q1CsNu9UQPEMQCdnoqBMZxYQoy2rp2
ipkrUWx2iRz3rxQYYuqbUxE/EqlOzMsDpDkteRF8Enw9UkpU6df4eGPg7EIZZkovUDvkG0MrOnPg
9a4TTCo1kn1mCn4Wtt1RQSiVzpuhR9UiA/h2FELxnmhzWv8rAwIGYnontDUL4dp64WXDESRODys/
6xriz456r5ESU6lJIz3X+On5bWDZsLfBK5gaA9rWgWbCV5tDD4wpM2k7bATYZGAcQ1RMsZrKZ+3H
OD5c/V1AN9UtCFOxYmuxeqQEXUXNCb3sZD1pUxkNCNuT/ubxF7j31OJon653OzCritr6DH50ISn+
PxiJwKaV5meI//JLyDrOYnBIst7+7FrDx/kElsQMdezROS/7+9Jcly04Rj6CoodKvnKtBFNIdRyr
9hNx75ApTo6Gcw3LJr+YWdypjMxAqELlB/81j0gBoEQtqkrCOaKk0W6a8wJa0zek8hmYSEkXgEep
S1jr0j9oTvfTbaA8dUBkbMTonEke0xq4T4ZzRnipoUlKB/rlE7XOmrqdbAgv2F8YU7WmsvwjehQy
5WfjVPi4YHFh9Zbn6W7kfo+/3Scsd4ea9SL+gefvH5BcRDArH/4cV3IRoWNfqkJkVf6SL64Dfs/7
nAFYN2FK8PqEJIM6TOlIsIhqhzU4QgGby+sIOTDA8olqua1r5Y+Slfy9b8UmuweJjcTpMHgsdhO+
JgRjhaQ9mFBv37+h9tudP36hOPVuV+Dlyp8FfFjh+Umkq73ic1Hm/H/w2DCTR2BoeLpJgq5wPOTl
laaB+4FPSDiUH0VaoHU2ba6gavwYp9OCQkRO1wirmXfatqI92ivuVH7Hul2gfecljsMy1WsECCYU
mK0OnFdxuiB7LD6E1+FWBlPNu+8d8o5SeYOL2wmtfRDFOR6gRX6mTH1mPzi+qQ12TW0i4cZJ6DeB
k1OqClud8KumyXFH8ckkYi4fOFli/s49yndGiU1wyrdp8OfbcqfOo/5QoXxjYhODQ+dAdIB5l0Jf
75SsMTUtS1+HLOEea3lnzW2Kd6exwsaUnYT/mt/xtdle+u9L59sNHCwbZrPuW1OOcjuTf+CGEW0P
spMLQTLVUCmEyxMpOh/snqXnAd0E0ldNjjvKa697a9Eq/vM22fT+ebhk2YBoiEfdzw5ERUTxUrMn
mTvca8PCdNliY5jnzqepbRk5GyisUPVtvAMkYHut6Dd9ETk/NwtUy57G8/i4iV7fDKUHa3evGIP0
4wSnseSsinxuoLPTL+L0bFsmhF6MYMCAfiVplQA+kqX+BhXFsj6/y8H2TwZmD+HORsxrQ4V5F8LV
DSBpg8cmljFjqYSrP/jsP2BluvBykKZvRgunQu6K0b+DxGEWd8bdvgBV597fNKZXGxhoSpu5LfDa
Yc42TBVXpz35R75vOB159nOlePZDx+AUApTYcHZ56769iFdHArEsbR0zBs1KvV2klFF0hWMPdunW
3LDfeXCrnJjG28zUT4wlq2tgfv9+FocknbFM0Kp6lITkx9rFxgJkAXHKSZTXPpS95q6lKLNL8pn5
ToJKVCQaTbvP6tZ4XrbN6WG1U6eSboFEtKjqUDgEnumCQswBX1rTQAQ+bto5fNHNU3t1fMM+KP1S
rqJryHzompO37oe4uYPFrs/tkRF96OS08h90YK9USrB8lg+4CaCC85Wovd5b+PXdrRffsW1Sn56X
842zraXaeP9Jvo0gULnrQaHkUcqJKLyJlGoOUltlNaPktpuEzCw3XKSPva4puwuNl4tip97C0O1i
Eyj+R7vBfJIc3Da3kkKsVmCwS/J06hOmDwwfX8M5La0vrCupbwU4d32+Yz3Dvm8MpHp/UFQF0AJc
B9HMXr8Kyv4QtL4ha79g/ov4ytr0SUvq4rmRSbSviIQd9cHfVCuatN4UKksC0JXrXQEu8KuNQaGq
GwdR/7+BLd7t3Eo0Vapa8qP6VTRIA8of+Hm9/5xFUc3+Ze1LS5ZTIo76/SRbAttptx/8+ueO2kc6
rZicIOPzpAL6YnzIfGy9Hh39xGytcHmrmuGSX6cLJertyZEd9MZpxLqfujwRYEooSNZESQhGMgF5
bZyKmauYaWVczepizrkH6/ppAFBkGSvgMqlhcMyB5L6/L9G/An1hW4XSLTmADTOETz1zOwN1Kux+
WBINZZYDyoIqSSp4CugDMU9nzZEPCEnCEjbuSQXspm83xEbHdM582YDznHQjuUwGArxddy1bdAXe
LwrI9SbhdL2gnrd+w65qNNBujOecqnFeARLpD/9Tog3osa6ohavR2G25XWbpeH0AVGRDwoSK6bbe
AAZLKDdY7oyrOoSmxE3+0ztObLdQbZBYEFXTJOuWyLIzm8un+IY17Ni+Dak7iw2CY7Mah7OyZJzO
DMHbqCjlIAwUd7P6qtMQkh/RzOg0HwJ7uUMNijawZKYfSS+oXPsU4YlmtDlCbd+5n7udbSF+BWci
2GzgwImZyYYeWRlC7dOuHQoL+nT6znGvfHHY+mP0r8YvLTgRqLjcwpKHTno6d6ysKCZlBhGBOEgO
ZjiCRjIP0Ch4kPHFyYHX455ZPAESo7R7R0iGXvVvpNKG/5Rp767TnY36t7RkO7Mp+8X5nhnRR7Ea
oXd3QXBhhbET9hhSQQd4zC9uqx8S9SXc+FxBBWBQ/QzHDtedZXmPRNL/wIjhlF1lWIxV2o0S5UsL
YUVJDCLErcyhSYiO67/NFaTqYouCL9EZuWqwMKxW+tV4OjlEr+jUkdmFdzTplJ34anXOQWL5lwzn
5RtNQVwQCWP/L9gcsB/ifgRJaEa44xT+oMC2X9ULpmNNlbPFUQf/303K6mB61F2/f9nWTBESZmCK
cnVAfpZZ92APFqHNjLrsGbYcnlFXvhLvYQeuAKIpJmS6TC8rnf2w8R14xmsx7hWezwU6fOI2MJ7l
kvFx14rBLUmwQi9owWlOIy6PUW0p+fuZPS7jL9J7/idYgBMg0jCLP8W4YAlyvu4eNx/x5vValu8R
ldrW+OUf7HDyHRpMCilOjtrubiWngEfU+G45XNb131Xj2yIPpCJmVWTAuRdw3p9nCrXz0xczsGBS
FvqErOOXY1itVs0yJzuy+pwFHCku3PH3gjoLcf9GUCtUZvAnj0BDCbfFR5buVcggCsqJJqlu8DMq
GaAUoMSH2diEH0yA448e1eG1VWVLB4yvBmoKAf0FMGdB9bo370OwIyvxkeUd8HTfObug+32xA5n0
32xLFYKtNe0vQrURNvox/78BbIRw3I+DQ39352tIRUdzrpq+8EYWRWEhsm3031iIcYbW8FZgf49y
EMmRoX1Orh0FKSHliKO8QzUObGgZYm+HEkkzVanpy1/vcn7nxNJPwdLY8ZYtMlLGxeQ+BHs+PPd8
hSGhOl5xRSa0gOuLHURxiudM0WxU9zK2QURhPb8m4h8bD9p7vUGD0PYBE9san25q7yRyxWja5f++
aagUrleEx68eBHC7W5ULsvocLVUnuAlAqS3/ZoIdt9gCeIw7KLbT5bj0ghdWUGjoP2nkdnV1nhVg
WJC8i+aIk9eciAEMxlIlcxudNwIn7avE1LFvhSKrHs6FR/bHjmK6fc8IV1FL6QM77rUvxyq7FNjt
Nh3z4MMlDAjIG/JFnYo9rHOq39MlNRzf8f/C3gloUs2fz9iIFj/wED9/o7FuX7G3B53YTFRI3+TG
qGuJZTRi+0pdh2fJR6HJKPBZzAMop4rUlyJyhC8FJiaIL+1ZA0JtHHF0jvFm8nPSKgcpurUHFnug
mZJgQ8FLMav9MxyLQGB0sCGLVqPvRROCZZ3ngJ7hgzkINOwR+M9EBRc5t4obzFQ3V3O1JlQ8Brua
bNlXfxNclPwLtX3C03a0MNqB2uxDfeQJ3u459w3VsTRQxGXC65RANcMI6LwECODerheA3L/Tqo3X
5C0LmJxlF5amYFb6o+3XWuiG1wuWH0jvHsneL3jF5IpdL54rBQ8Y+cBqRwXzxWspZ7LpnCzgwDJD
BX4KbyjX5jjEP3BB0jGIxU797Ucr3Kk4iqZKTy65qyBDQpT1JGbFzuLrTPFh0zB14JNQzCTDzBsT
T/wP4/mUfokH6oUPTRTXZX/KYRPjbDHQ3Iee4UV25JGjZGAA8QVRFcmXNSHbNebltxTOh+52vR0m
lCAnSjYsAHByK4heTrZSAGOdkx7VUeoMjGnLFMEksJPyt5aVljqQnNSkcoJg1BhF6nBNabp61tzP
Gm7ivFYShS9Xbc8VctDwRdxSSbAYeLVvptXG7GLV761TPMx9xIKEQdRe/vcwIPA7EsiuZ/8rYhYh
9nysdFUt2GepU5rjVfvwxi2u3N9wgABg66Ae2LNHgYd39Av/skggXrkEE4yqPDu/ADVKiDOxttk5
xnu3GbHrq0FyEqy3Ao8XIQRWSLRrOi3vgXpmAgoTCPV7eZxZN1vNb9OUkvZGs/aj1+yot+vhd7Dt
U4BHr+USnNuiR1ZoM4toliefyi/0QGMgAZnPOOQrY+oQjUmRiT/To4Am+YTL4LWkekQYnL1nLNUM
E2CLHaQr819RRRKiYFUraGa8Yz7nZlAOUftN43+ifQzQFtGuD0BN/t//ct19XP8BjI1LKAwRvuF5
i9p836IgRfCIJ6syQYyb1dgReoPJMIra8FYvi9R12h80MqkEtViynvz3vSHrfeK1Jf4rKZmrCl7Z
J1OShp28TItYoY+Gce4HUD7h1c6fPr0Oy0JHbEovKN/w3WLqpP0aLwtmbnQKBW4MPbEBS9yjZIO5
eSg7tby3zevoq/cnba8rmACK0EtbkBZE0dd8y0CiPRXpvtnOuC4EzAj+mtB6YvdcqS2QXYjTcd/e
xLnqZmsz5Ka7Ko2X81/94bXMEw1vhxisV7RpJ7WzyI26JM1Tt3QcBgN/0mPYM0bZWsqT0cwzk3Hw
2WlM75gbMNk0RJ9XoHT4+GlPTwzFgsFcNeMwTBhF6bYvm/i5My7z/MNci3Mm2sWxRS2z9CDDn/JX
OWUiLjeVoCmVwrkKXtbvZDnLvqYmNdHlBZUXj86LGZz9P/BP2CY16oP13EV21zZMrAIIaBIf8Ffh
Ac80kOM0LAdZphHJfmwCzdKfQxzwzLNlZMima9QJKBEaehnMp3IcNhLI6hhs72VDBMaazlu528qZ
3AjyiEeeb3UcWA7Y9dmYoHstorA28UFMixlOe4esw9S+fnbG7HMlMrS0CtzifyHq6rGQ4BcB4vDl
M7d7mtMfmm4yTFKEc11JumGJPaIsz39vMqWKyDce9DmcC5bs0H7bF0JunZLgEGybtkf9tjZJVoHl
6CKgSUdANTFw7OWIxp0m8tsyo+dSMp29hpKI38NExeAHJpcwZO73ucP3tqgAYukZbtt8ho2EYrbu
CsH7yX1dHjqW2eGGziHZk4QnFi1vTnOZlHtR2Py7y40iA3AMGuLqzatziKB5939rNwtY7FpMIqkg
20kVVvFv0tDUHeOn8yQs+cHU/l9JU9bypq9bYICev5Bu3y/uYD4wanBEdLa0h/bRe+PEQK+H2ztb
6CentLFCnWTM2hVLuhoZTJJKPHHWKVlIkXjSa4+bQydZ59rE5wqvOuuR+dmK7lIUAoN5+DUaKEjy
nYyC9V4xTDzIuNvkHKPnzM9E+RPN3oySbQpiNvyuMD9Jwz7p48AJaFmwsEQLsJAS620E4cWmIcJd
nZNrFCAPB50odhZTUPtJVgCm8jQ6L65Tz6YnkXLY43mu17nSzTVoEyodm2YANk3BBr1UiHG9MSx+
VXaMpdB0aCbe5xXYaynmaXJPA8NCt47VW6am6nL58HJL3/UnNZZdhOyGzblBfHdsPLHVpnamf/tC
6T6+ZFqbqzFW/558+pB4mU3PUXyGP1msiAg10vRU1jmH08syal21BZSqE5ndbe1h6JUSF2T29u/0
dI0fi+ZsglFVTNlHz9zJUwYNUYGbmYEpgYcF2yfbUShWt+IAOfbh81+RIBgn3gWP/W7YdfFDiWdg
kpw4ldVYjG7pF0M3PZdK5uGmFFt53hnhCS40CLl9turuS30lUO009GnkFl2RLv3sZj9szAvWkMZE
0mMXGX0S5+PXONZeriKrqTcIm1ebhyZK4iElkQ9YjN6iJboI2FTSxQVLnI2xO/VJ7sdaZciB9zAp
jYF3OLkYojYWy55pSE0ktGh8IfB9WclhuUkKpwOgP6iewICQhv9rqMQkQaNwmIPxCRJ7g48KU+7+
xoSOc/jjK2pFU9QFxYDdVxVqKIS8HrDcDVblI6dO901qMic0umuh08xZXt83G5wUz4VuDTTMcP0O
pLKrM8QmSIZ2mFrk7OdlHEqLOTuXG6LDQAVFP8NHCTPaXn81jn7LnewqSNrlOE+HeoFm1Hst2GL8
YBZ+dHFT6E4jKrCCIQNKcB6bBl5N6Z+p40mVTvWt+DKD5OX4h3U++w79s3pJ/ALGe9ByG5gxqFT/
zUj7eF4/h08vZoxi5vfZMoem1pPNHXF+q5nS7SZ7jK8U48Fss7dxYzv8ePic2uZyOgmqpN3CWHk1
zEUBrbsyBcQu0N+DbfYdlJKsP/H1orHj3OhMGCmsMJtqxMaJzdGY7wf89p1/+s/lfcaVgx/3MT1S
DkYUCVTOKoqjqKeOQznPbA2X89Db2BOq39FVqKe0ckW3E3alGu4x0ciTpMg0qCbQUreub6IyIgL6
VZXa6GMreQl3T6eDyAO+mdnGIQExcTehpwbm9yzRM3yeOiV9yIyhYtm+HiL4kE2WeBu9MfE7YODx
A9oizRRRUH3QO5ZO78m43WOHXNAae8HODZoHX8Ef6YvuPhq661+6eXA4oIGA+9LRvoAksQ22ledB
uA86jpUzqbZOBPicJsbl+QMbDpD14fDRBMHm8jtZrMmzgi5+bxmUmAVSTsNIJnUwRL3+cba0JkTK
niCHq8sB/T5/OCxmmsCkcUa+Ci8hSa5sVmouYl6+x1/N+JcnlbwdZBfNXdZCIWvGaqa5XMDNx6QX
6IoUZ/+sKLRXxNQbS/GCbbimMNFaoZBQ51wbGPFbGjdXN7edxXtmFB4Lu3uupsm0kiHZCef0zO4R
oJJNho6GAMg7Q8KKVQubEQV7ezTuEEdZLm8qdNU0Lc4ndUC/OC/XRA+mkin/lIzoNx0pHj2DFzTQ
jmtfpJ9jVtkeiQq/nYEtuBNC0rFUa0JWrG+mA8K+dlSt4yfU+JzOhApUK8XmpAvduBhoTTHIQkHH
yhpFCcr4LRnUZMMT7QhNtRIA1kdF3F5aPbjpW02INEIi/UNQL6FUAkkfX7/AXhgPRu0SMizoHUPY
jauWy1kMpyMU48DgwpsVyfR8BwJ0m9TS2dzzTbfxFFXOjweH7K9AoJhP2wZqLHkaZYNMO3HZ2bx7
7gZ5TAY1pQb1Eyi1P+QTD9Kt+dzbo+EP8dkxay5yTi/6Yhi7e60/3SUI3RvhC7icwcTiqNboyej3
dFkwwKqhk4CJD8J2pB5pAGDz4aOW8Jrbs9xRPc1wLr0hzdGDRCD/FC8F2KnkIMW0/js06OKhdqe8
rrfLhP1NXWaUnenk1ydRbPNy53BL42A0xgluONGzUa4dtgO0thfXc3RZH3zFgsLG48NQAs784dL1
LWB/GNLJ+DoQWphQc8e/CQqbJYsl/TuObH8Pf6+127chxTr5C5KBq8mAnDBrESrTwfPfp900IV5b
rQEEXFEUOxUg7ZS9Zy09opchE8sogGIKctA36igPKHWGBeaMhuy/SdtGr9HTpiJpmMF6Owig5XtQ
x/kHVvxX0dJEemuA+Z9XwzuEC0gnZgEchAcr0ZHI/Vrh78u5sunsZ4HK+Xd98F6otrF+3nPsfOey
ZJyv9KZSO7gqQI81fpQmAFKmefwMNGyCmitKudH4RM7+hOqZW41pd1Wjr/A0ucUH+xvvk21WhRki
WGn4eCkeHfdMuzvGNloLRTGMfayPhBNkcVXjadVObUWpdkQ8G2awoRyjF6IsIDVVi3x8WBv+AqKS
+lhWYqh9FLM0VvrzJuYK1i18PZq2tT+MHv7AdyzBmAs0lPgoFh0m2BabnVt7r5fOn4pZNPXaRvYo
nuJMiRJ32ixK1vRgQ8HzFqnmyNefLk+W40spUvV/HqdUF2XElTSHOVbWRhvtmrGJ/hX/V0LTIuBX
987a2QZttjbfMLFjTz7z/UhYIclswJ1xBWIFI20eIcB+/2XafEYbut7cSoy9XE5z/WOx84WK9Wx+
65wpoLp/n7bfCAb/Jx5qdR68oS7qNtraHLdXSCYqS9lH/oVvalgydSLcc/J8R+V93h1RyRCNmRuk
9dKUSVK1tYjgTagfy9sXstklOtu8Nfk/7UwGlqUKjzaIckOWsR0vzti80ESnXi43eqKoBmX2ZHy3
7MogIFVoOLoxIrWlj4PTiErUgk3DLtXTQxzOikFlpMwGqYVIh+jEY9F3SGfpFkjUi9rut7vozlLb
7XgF1Ru9twL6l5bZ/Z4xOpJIf7WAyWOOeVodp/qqMNBQVVOhPOf2u2RjVEta4f/wz+FlDhOr4ut6
IIWGDJr9MgZ1CYzIi1m8wYTORjwql4u4t3+PfIO1mYHqQeeKTZ/nvwm4U6Qn0vpUcPWLTdjbFadB
vGzpdF0dnFvRFwLDZDd7qsYB9gt3Ev+IOi2MwqsOBsp5h011D6VE2p/M5KZVnieGD76SvTn84hWl
DE5PHUEL6rgeOUYeZM5tYzpQha9lg3wc9LZDfkWdNTwDj+kwmGmlBYm6eBgYwxLVRctgOPoO46NP
cY73fcKCzvxdvsZC7GI9TzMdEA6hQDizNjoO+6J1Am1q1lLWMct1WyyNvrAeAxvXk8X+SvFS4wxJ
Kle8fb+wokYBPB0fryxebX4mxyZYAeUyxixygdnVcXUvlqs1JKLOj1sa+2HoooHCMegF0a0Lfy1y
fsIuAVDni7QRqpJku56rX8TVHoxthPkTcaihgspE1pxLvaikEIKDxHnDRcUKsaeFiTqOOa0EQhUY
VvfeDntoUGFbvSMc8bieNIMQuO5FbkVOVwfYXDbbTgPDm7RFuDoJwC5ii3VoHEYIVFPoCABgkv0X
7ON1w86mWjwZ90bBiAeAi/GimRMlBsX4q8jcjV3pUVYxNeSvJznSB0A8wD/GL8pZ6CZgR93IgFZ0
tArnUzaJFQZD8MkKATxzIvuJCvYH3eL1/zMWXzKSvuwy9UID7HYKGAbxqgi9h2fPX6z9ln2qBHTs
sVhbM1qKpHRDW+zMuQZOmc5cDnqqYlIZ38zJrVDEU5Rp94QEp3KjqcYZWAqGGo2hu201iSgNS7lz
1rM5UMyCLv7vfIqma/qbyidhxev73N5VRufL7U1AzjA1ljUktkc5OPZPjYmTeOhXtZzDrSQqDHji
ivwL8a/Q6iMJ95Phq3jZ3ZdqUOr/1r1g+fE4n022obtSBZsoimSx259jHubQJAOky4/a2xllJTbY
JCwTAThhCcJRXotjvEgdllb6bIvieF3QT1rYAQtx03Ji6qVFT2riBjInyDtyfl5jh4ypXwNMQazB
hgJkoe2+Ob2B4Vlq/s4fbOGTIt2f9oqGrjFGXgC6cQ7UlvxE7D8MpaWesWE90sAHwxu9iYvOxUw9
EhMfB/tp57AAY30wiLr4LRXcJR7TGa3fn8H3EUODtkoXt7GS8JjlrnvL2Z75FEUTIl+CYieqbSSG
5umJ6M7tAGmO3JHUbJ/+Gfbket9+d3c8eoFsNcP3ROCh5esBMi9LW+fAAGc6m+IxHUwOoV1C7TO4
KO8YZgE1Mc91uuJW2l4l6tengxh7SoWiWY/AERWHrVbyOiveeAVUt09+S397g/P7tiqpyjAwIiOg
VqE0R/Q4qeXjS0UOuXzTu/EcDB/7pZ+4oRhRALr/zcM3iPvXAVlCkMSgOre9TejnAKbRb/02Fao3
KZrqsc+zJjjNJMtwfKaiIga1Zgh9h/rKYsk77qJgAxdlSVAXhxhMYwLUV8b5bSTMjG1jonhLYRSb
Kh5m3uzg/jEOIG5Pvt4vWlcLcvHmMI9vr2vCw9IghGgRi0z9A+mkjgs/fPXONayiH50w5JkS68o+
S+nLkuOmSQeMH6zN3KAkWgX1b777hG5wWV0J+wrdjsRWmwiLhKGF2gxfAvmrOrDOBtbBHgYCdQeE
sVuvh/NDRJ8tBzLozmGGSCiDz+ftKnSHKRJ33kFv2rd4b4THAswFX0x1Sc0zHNUnf3oV+0xTcz9q
HjDZhVTTvJ3BSsUE+tqYPH2uQHO0MAMRw74emGcdUqWaZNIbodMiidfjnPDBFqZ0EmPuUxyiW0fG
Dfy4tQffDk1b2eAmJHyFC44NkkoYDSzbViZAts6w9dqx3CwJx8EA15Kwaw0VgzHRzKvGNfN7UD5c
5NPdHeAtRzd/AFwkh6G+vddIGf01WzrxcAhZG8nyzdiL1XG/kYTJp2R80yFOphJjV9J4sXHh9fbL
9+eFBph7JrNT9PbcWCKdDmQrKEipjoSwXE+U1rxhlxXUfaLW8gLM8t8Y8NBN0Qr5PNicyP7wIajh
ofalAiQaQoUEjdUM0lcVnOmHDXMoZ7p+dXy74QEHmtCsCU3yn1cCEv1B53WzR5zIiUVZPNSJsIlA
ZcH0Ch3SK9FcMDFSNY72PkcSYEZWMbCv19jdj7nufDnVBvKbs4fnzBjVVNWuEP55dk/+ZP5ikU7G
VDHjrhx30COHj9gdbJFtR8qPxCg5VCkMSSpvwjt7urKZNeDmYUgOWuVXsi7y8EwheJVK/33Tbsr+
XNI9LXtXWXxNEdJHy04M6UMMDobOK4km+Zfle/9R9SgruyYY8QiIBvoz9d5fPIe/Q9KF3PghnxQR
8/4AMoFjxtw39e7z9IX0cw7WejAtDrgzglohGxibgOpwEQSsZ4dURFWZGYlIUA67MnbwisOx4SJ/
WQPVX4UpekxxjXJfQ2NUzgMsel7CrEDffYaL2vHJ/eDihmwdVUNbS2Z149pyS6LuHObU5+5SLx6D
x10tvKa1P6OMRc9bO4h+YyZdt9bpOIKULyfQ63kpQIXtEdQeUxikmmGCnsJNRPRUmQgZ+MUxNiRv
uhngaAtcbHCpoMXewNw+CcWzh2LuCuKBexOmb33S11bSfftBEAiNL75fejNZvr7lHRTSES5k1Gkn
tDaMh11E85Y45SuFyvopDSPlEPbAPhVXedP3iFEHpKdWOaZtTbfsBqJmSbIo1GR2rlCbGABnRlZp
/dt4nzIyKvZRJ4A2qv5neUG/Cknid3/mmn2aSgLhcLqH/1r95qgYgEH+EZ/lzZ0lyLJ7dhRroyCi
Wsvkuh9MkAIKRL0ejtqfE0UVFZN2Ufde7k8VIeiJQzDr8K/sxOZRFDVJpcAWrEM+4JhvUUfEkS28
qmSN1EdR9hEvGwEstNiw/ifTlWN3jnHCE5hyihWiOsRvGGrYNI5aeBZWydNXSBd7ElUYRMH4FDoW
qlIHJ9fbbHqn04aZ3kIUVgzO+CLPKqgWRE1NpBTvMD4f6kchdv2Bl3+vZny/Sy8t0p7Ar5ppXPhG
4HEibFBEPuG9UWv0TU0nanAnysrqYNTTNwIQrKR9fRthuHhv/n/y6W2VeE087jr/nsLNiJ1Ue0KV
EvC3+fJKPUfLLXrvoGeds7ysc6WCJX/UWm4cA5Blz1L1/kmdyi6lR1mUdG0BXo8+OjfCvbr+OGyt
7OFw8nyfvv4d2bovaiMvZCxDhUR84UFa2kjuauM5ryRT/7/YPYPQOo2rb9DxhnF2U1YQdAoXBBqN
s4HqClcGshoRLbregbEhxhK5n29kDzQHFN8wZdcRM3iJKIoXiFH+4geJpaKpTOaBhyNAbfrgRog0
V/yFtuqjwlOBhR9pYyOcXQPv0YVKoUcXQecLrta51RNTaRojTj6bko6EvEbi9QseKB2MEzvuXCVI
jBm5fRP6hDQaP6bmOmYrhIse0lfYa1cqgL7+pM5hrF7S0BGTyUZuqMfT7WYlZ/DLdG0KhifoJYYx
KtNUnaDcv9Sx+LWPOs7FF6Sr2hL7eRRIjq08dSnBOMfGKzNpCwsKS73aeQnRLQc53waQPDug+Hxk
fsX6aEWrstX7IBoaOD+E02JDf4sULSB5S2fKpa4doB4JlEaNspOEOWEQg+YliksGzfhzDNb6rwx1
Q3aeS3pElxpphPa8yDXq1N1W5bJqKtro/rt/TRDgvxs+WuRNSRLQORMfIWluHAmhySrCs+dIVjz/
zCuDJDos0nYHxpihY87EfBlH8IRXWHkpQZz+InaWscDYpaeK5Ei+HFU1dfLsbPhJ1nZ6PR1u72wE
3RdZWP1RJeqaNxQzTqtkY83kj8VRwFtKUlidWUB78CJSiegXDL0qzBTViUd2n/1OtAb4cdYY03Sa
CPQrGg1FZq6u6o19CRC8KrURglQ77KdEj6u06nyVPlLz3eN9M+6WnswdHq0woD3pSbbE4+710gS/
aDsADUFgwp3u1XcT9yrpcugzs041Cx6rWEVnBp3LcMMcfrvgrUa4/FiE60WN+Frw99lhBgPzqmwL
dsrpJv3AyADurYwT/idYzg06HS3B+Y2vMqHpocIZWC6KFvMDvAoTc0/vXPvQ+j8qgntoN1kKQRil
JVA5uN8l8BTVPVIOedB7bL6xrZXSRuUu+SGl04+7+3lOHu1ERTwsymm1RzHw0z/gbbPwZJfVNedR
WqUBqTz4xS9ysJfIVIkf0GzerPWOQ4mbEL0/nT942s/+21FFtzn5Nxsex3xMYpDT5FLW8dSArohH
gMYPLw07817j7OXb20OAuHiJf227gvmI0zadFoASr7xfmNQRat/Yan7aMW6Cb3VjKEBO1gKFpDXw
DMvLD4rIQAiLC88UL946KkjutEFLkbZbAhEgkbpOed5/Lvqx3YTvmFh/HmcVhgCrIuzExGmvaXzm
8+HgMrU6wQVJNt282h7nmEx1rfVtsALpvfWGgm8hCcQ55yl/fkThtXn87HHRMZEp1Ay89ZRJ2tnV
5Nc38VCLbqLuyhyNg3ebHQqRW1t7TYAkXHP8Vsv042wVZ+tS19Um+pHYZ1EvUksPNqZwA7zMzM8S
i7hEGK5jQa8C+dfqs9QzvBKEcyHcLPsYfh7V3Ge/wEwU7PK8XrWVWl8QDWykRsnYCIH2boQm7KRk
UwPe3hxKhGUa3qlwhwzaqKaDHJE8nU7MVKGAOmmMv8YKL76sGL4wq7LGetSXWYpW0KV6FMvonWtF
55v9va76NFe6/DTrLg/WOl9gDKuKptkTX2UcaqWMxdg1YzsP33r2htXGpKKRPGBU6XyjbJwyWgQV
hJKMGEdo9rY2yBIFVuArp4wwtvDGR0gvF980+jtNKvbbNmRI9pWxxm/n6gUpqzoXPeJEXwXDSbMO
31IOyshiKquemDD8D3+isvZT2ZkE2NEDfEqfsGqtHc/4NAl9FAkSZoIqaAWIFkIy++pZd+7C4+vf
KvTqdXRxjkiGaN5tS9c5N5k7V3va+04sL3pkfI16C82qckivqMb97rTvm/ywIfXi1ekd4TNUYGKQ
YwzfWjrvPK7O2PjFjQ+jp3W9lOifQwLCAKjTd2Qo+YPE62Zhall6BNoaUCyqZAnqjuf0D4Jq5IdG
D6jKfIp+7qp9uHQjk1xyXDcUyrUjQOhT7JuPpODBg0jUxzC2nocO9xY+L2qehS/kYZPTlW1Q+8xy
lJX2RdSVapefOPskaCG1UUUammw48k/APZxBHxWXQfRW77Go73ee/50G/YBYqNHw4JKWlaKzCUpS
BdvauDplNGF7hAijsZnK46DDyV+RYjk0juRuaALvqB5ujrfoUOqR2qVeTKkqJNzZotiEyU2N/KSt
ITFnsEllp/rTsctjdV89uCEyUeNmJgLlVRDLG59YDYL3iFnJE7akDSl6JDPOulXGbiY/LQt2xys/
fa0Tn9FRMrfKZwq7x3UuC7go6hr+pJfx5oA33tS9xX4uiDwpmLTzFOjOy7cHHid79RPAAl7bxCoF
cEPWebVETWTa4JvhLdal4GmQTuBYgQU9jD+Y9B+itSG9jKPgumh6Oy0djuJH3CSa4wJFzNm9hoLy
fZY/ML9ObUmR9ViVXK/Qqy+Z4r9BqNOY3gbndlrf2bbWiBWQfJEnhqCWZN80azen4PybZQk8bs7K
SgWHt/lPKctkF99HgsT+im14D3ZYwDRiPtJaCud7PqNDhXHnl360Tol5JyJnoNgD0AIDwrbk82FH
h+OJbryqOLGIwyFpozHNlw1/EKwAPbYSKKpzUC0n5Zy6byxw0TJUh5lyYtiCLH1nwCEodRB3fjYt
S/mW8ncSJ/yvzNQGRJEN+OqTFtM0PLU89om6l8tGWe/+BooMl5+eV3X8WMiyC38HRR9wOyy6Qh/M
vtUxcDiYG2Z9PUAGOG8WwT/DU3HjKEnDWwVJr/+Xw6Nk6oMtHGk8TL8muIhz3EHzu9j4BgzJUare
5qeWE4odba5lb0lhzaLE/oZFrc2OQVgwyleO7Xvf4CePuDuRSkE6N7hEgvS/XLpzWQ1OETV0QAwa
D/oYrXClEFY7KWRvkPPRVUIoPAIpmIOL03R+5s+UDorDnITEkDVncLk8AhMxPfT7iR+A/B61i35r
sI2/IIkF9AbIcBMBfWTUoEbO+V1eMoCDh2X/UL/LwGh+j+/wPprLfDkqTbKWcyN7ZSUxTLEsTCT+
FZi2sUbIR8TXNHjvZbLeJBVZO+ZsRJyd5ZPDYqS6hQryXdRdM5KAX+8hWZNEUN9RN4KgS44UXee4
EwKMIQIFeEr4MoU61y+3rsuJYa+E03XFPfXa1zr8SCLInsAwmUQsgcmD0762e89ROOYub6w8QW38
Iiz7bZvz/ugUBMqBLQhhwopxbJZemq3CNklfguPJcfbt3OevSF8LkZDON4HgZJCHcE9JuRAV8r/2
jRwNQhy4Vknlv1WfCuTbJlka6wG27zQmkn2YFPLrRjivDXSH0v95LEBvRs/QR7jh+TKdx15b+z/c
bT1BbNvs1E7LqzAyzfI6JtG9/lga/zapIDo0Vp41pnuWKMiS5YOhs5nqxwYGOOVcP1zWbFWKFDnJ
qOaPMW9fb5iOJosvK8x++LvpRHl2C4wkkJ0cT22malhR9D4WK9o4D4+zbiELGARe4uX6JEhd8HtP
5iEeY2bsIEYGilHtWbKU+QU1UoWgf1xseI1BmCviMk8B8n/oeP4t6T4CHzBBLhOjEK3qiz3ZLMND
ECHSvTLU7+Zaa1NSsqDHys4UH0/l3FiNi1qmDPw1z8qWG1WoYyxcRf+fJ26tUoyPUhFftAOPcPLN
oNPtO1SNlr7rISoraCDlH+pzyecJsQo/4Jk+l20ndVDo5Of+AUBIYCvEOT6IWJgwokF9fedg6bA7
1odXMZE+VoBxpqGHTbGuXehIEJpmULRZcDdTRn3fdm0EZArJ6wgJwlX1m4HQL8SpQnHvcygZgOne
4xlk+Fszpkb8aq6XPAp93Rk3CXeppZH+Gzu5tRyqc5QtWOLfELmPT2jfyO58Ya/4hq2Fyn7gzwGO
XX8szf42R4RBLeIV4/qs3o5KDiaBx36lJaEMlN0/sZAQe34RDREM0WMIx2fLeHLYVeKBkgAAGQJc
V8Mdh7PSY0CrQYOqkVHq/3Ip9LD2woSYiInOGNV0WRFfkBYcBAqpl5mRig8g2ZIH/hDEM6O6NZJp
DtsfIxgEfRqK7UTIv6rcEgsRFCIoMN0urzIxvh6n3jNtl5SumZzYBCT2vM0yWQdmeXEYC34HUCdU
RiZTHmlBWGREdybtLpI2FSdm1uFEnVi5E0tmhNxZBRSEVInu+F6RWUF4bF4Lq9R+yZMYxO8ll1Vg
EsuhbV7Y7zmx2i/Xo3ieoJnhnOPqWr2RepTe/mQ9bOfuAY3EUYjaJOec8ONkrYgHM7iVlQ6kS5Xx
W16mWpAuc85rzgbAieue8bDzM0NHJ8ST27Yds6edTA949A5AChnRYttdxxPFqJ1nubA94RLcr0hF
w/RTaF+A62JGaHfM1XeYLvhaK4/dRCQlfPPq2QrZLdB2Z1oUbGy/cU/tpXhwS8XUTosudorcKVB5
yA6LUOVMCGCi9UZtb12gSszcxUkCjMogvxx8uF+q21m01T7ye3qG/rYc6LpQRUkAVw2DhcPF/MkH
c+TKh+HrUnzHRZtBcfN+c9hb7iAMMS03NPTuzXpAyG6uKrAlyu7h1QKaTtK7Xb9BbyMQbumv+mTY
NDI7oPs/anQinVnpQ8TggsVuzemry5jnocWInTESYvnKL4PjgX/V6dsrKEkh/B+h/XYAJ2pZ8nOd
gK7dSJwNQx3IdmNJR5BFDy8EBs0i0JJdGV2RJDzO9PUSMCL/J0B5Bf+KN64ayDH1ADJf6P+OX2Jf
HDdvQRwuAQFtBbilyx3+2g3YHU9xTFljZDhnfTz2b6ni5On26NIxuXqwMhR/4UvHGpwstxw1cw1t
9j1TFsNSEplDR2bNLMrYzYZDdgmVa5r/bcX6FZ4j8lSbYvik+bIZlA2DTQe6GqSXqCtztoM75XcQ
RUBwvuFmb+nDW/fJLUovqrAQvJ4VfbZHtSFHtNANzQHT5vj7/O3J+5VHQ29HymB7Ffgp5rtAvJIF
ItenZePhnnhpsFjgSBGSgEVAaOJ1fhoyhBg9uWfHMYV5Qb6ivc23k7rqO5YfBgNx6qihl7ST6SZ7
X2r/pIC6rpC8NS6XhKj3JC0y87R9IDR/9kF3aW5RaoKd3qTIQ6ClxuVCjOYAzQuXtV6rWosWRIpF
uPROjn3TywYlRgtMwbs4lfMhVCHWRLRIcyJDsva7m2kNjUrZkck6GjGCqgl+HN/ZRQeydRRypx/f
TKUh5qn6gcAF0yE8qXJBdaemXv/ZSxJzUpMdU8uHg+2YWmKv6oguDSOUyVYnw9LalfreltQxlSoZ
EmYR73/OJbmLHV74qw+IdRqQN86k2ywvfp044Zdzt93iGPf45rXMSMIbC/Ts8O06uLf2ax8oezMc
k6YHWyNCecH68BiYCcr/Tax4dSumzX+MnwYhsZs2jjkfwLAp50YOEhjpokR8L7gz3dVJYYktOMA2
p0A8sH1A5uiuqmRgJxHrpEXDmxPafk1e3NN/B0KZT9FLI3HqzbNQ6WPKO4WY500hMYj8RkmI/2c4
ylVawMb1finlCZU2LKeu+gKfIVctSL8UL+ogjErxpHOuqOA3yGz800HvKNYk92/kM7jtaTaPIXNC
tlOBRLqIK0DoQCsn7qHCaW9Y+ye3WustWzOmOK7Z5eGdLtGZ+CNES9pHF4LD+B8ml5H5+JnNig68
nPuJqPH4l2snnYcttMS/iuyBh/tulReLmuXz0yUG60cpSIXupKhkW1jW5Z+rcU0LLIhPdCZSKZvD
S4iI4a4dcPA1ZxZrTa0mN/xXMoN3CLFsTBRXAqBmTX1FG5sHJr+Xm3A+o4zFAB9iPIRMp/3HPhY3
PyP70qEzPLDsZ1wMv0YHhxNTtyvWcsPF+k5P3vw7jioxIbpwiczBqVEmO8Zidl+M4zPQYY5KBfZG
huVcbUcKg/CqSky/JVSKx/+kjoiwOFcuuG7GpmvRFerzBbGL2ZqxNSntufLDGSqDA0luTa4j3jlH
e3RUUADJ2/qKCmP1CqpDdLd46ESjnEU9aOzDCcyz2YBTvE86gPgw+NoxvIyA1C1Q0mH1ikDvYe4r
JxfN9b+EC6xxwew21SKL0EPthvLsxdvjggK9L59tllgwpKqnPT1vJLkG1CIrKAI+tIAmUrAe5kjb
Ht/8kmMq2NVf6X3taHIQ7/7sZSFGIRzuAQ6BgpWmR3IWyI6+4AnxHhyvt93t/fCFOCo/SZ0HSjQp
2p0IfUF/AbtxgEHhtr0f+lUgvO8TGBNTkn29454mTefIYWce9yKOI4Z4M7b/ht1RLZ1yaoM55gcm
Imm1h3YFderFfRhQCSmJdZw+qbebjROM7V1yibIdbSwMGzDXdD0xysEhHlK6P/KeDZDGL4LQG4dB
Rl0oDIcAS9UqRTF8IbEuDlgMzXCN+Q9HHBMz44XXi3jQOhoLy2G6yw6jcfExzr0jWuXbCebAADH8
PJiW38BR448mXIGa1rmu3YJYwyH1ktxmuZz+lL284zwVCAAMP6kyo6lAvo7vvzh6TiGwYE3yxfhC
d804MbbJaGpajKFAgkfNaThcIDsMYHu2Imki8QNaI/QvlJIs8NohUYQRsWxoKwVfJjwlwK3zAoug
GYU9IvSlm06gshbNEDpESDQMCKVQ2l40dwLLSZgRC7AbKcuzE4fa/29qMgLCb2OP00GN4EIJxC6c
oBrBME3sGJm68fPeqr3gLgJL/m6jZwmdmAXYG4GpWOePSLHYBHsAg2cgIWilYrq0F8weQ3zJwq2d
m2iIlgay+0/XdI7pQ18hKNXAnLziCkspf6JOWGxvusQcoEh6DwNh9twqu5LauzZhsL4f7Pdts/jv
j1POj+ehNy3hoigAHMeSO+ICa957+Z3OMOmcM6lUERB047wh92/OzWwN/LJmqQ9CGIaZqJiwjveW
NX05KBCWdHipVtP7qyADUeD+X0jInF31Ktcmd9ydtI48wZemnq/U4eL5xYcaKrIats6q4EMKVJQ1
5ptyJ1tPS2PqebtLNn6fdv7WspSNdU1rX7A9OfDpKwxq12cwk5ldqmozHlID2wU9sdm69CrMDowM
J3OfGal6I3/OFJc7YP/QviMq2Utnh3tCggciMx0eop53UDMI/ImgyuAGGgdGq8GbLczL2xIRCnxa
aGvNnhK/BqayRyIooV+4Z9AMrOkokLLr2zkyvjidWeD8H1pgJmxT5RGiUw9/BuZtej2FxEofCL8x
iUwCHXiwMmSN2hgiwN+ZDOTSzyFHf+JZoHqj3kGfEzD0aWytEuMsOlPfFn/Aa55avHIIYPyWADMv
wIHwaLuRXO0dirgPTCsPBgV+EClhiP48u5CsBj3ZQ8dTFfv4pXbv0tr26AL+wbl7zy038s6iGiq8
lf5b118wwETNG8mwSk8hnbTEd4awUIU0k8BAMpRoMCbbmwBKLjdpBFhAZXSkV/k2cbAwT+Bm/Nch
gqTSJ28ahbdzbjWwdETuBU+RmHq7VushvFk/cVhyzTJUX68NfQKGOOcIv+6FpCK16gm6ng2Qk3da
L4Z/Tqoh2gc3tCCm6dBNEBHEt0XGDgQ8xIGUl5bOr2odwQZCN3fkKhWXSmS5NgVo14RYDoVxwBLY
QBOoR4SqPVrE26OZwLjm4dnaRS9OWNAquZBENki7HQHl8Z+rwrRjAyPiLKIGqHcBPBpvi4V+URc7
9t6mkDyQESFBOOYckR0o7Poz1y7No/2CqsN2kZIB37d5SBk07XuIDP6YGt7hCNmdFpVfkfLaA4M3
efvmLijDJXXK9xpNCk80RT9zFoECncf+pdz1AeGuixOb0eMUu3rppzQ2gcC1oFIhJxrOwEDpqb1s
25wb1Z0PIIJO9/J9f6XQ+cfx2UrlR3qqBpTVhMj0BL/rs0a9vzXSu+/d7nCiyOM2RpQy1FNQeQSM
+5WYSzIIbe/0zJDXRGigLWIzGC+DoHVfcHxejqIYFBnznjFJcItwLEFxtUyLBU9PD9Q8hF5lfa1k
tntifQZbl0wi4bv7TT7VlR1mZiBI4zV7GRYECo+K9vAgZKaOAyn5P5bADqfJ3COuSrCTcka0vafw
NIbCi9HLJijuliZMwnPrjDVaWiw1+cvLNIumJwf49Dp2jm/S767RURab4t9vUihZ/erWGh0rMUyC
cZ1BJpweNdW04G5cTInmerk1VOJG994LHUQNhLdRcIFpMrKjTNYzv7mf7J3z27FY+q7KLBCNODXn
XgVaYjOPDsX31ql+PHttDH4v17lbytnKnc7D/tuSOVXkJBkjNzMhJXoyPyOPvJQlB6moJSiRki91
dJuLdBWfWTuRfOjclSdJO6vyQf2juAYQr9bCXxLgdXabxIEf8Uo5DK6w0/17XQ8D+Zfm85+IcJXA
BPkxipojv3/HI3FQVQNLDj2hVnmRaLqMutZZgq2l324BKpGqckafYoT0AI6CuZ1PQj9O/smLDE3K
hQE1NHlBV09XupFcAiA8Kp5uctcYaOwXfeqnjUI09UQMn1hmX0gXkTItXCJKDVv6CaOJDuw9eD23
2yii9PGfXkhLHfsmqvljthq9eqH8kJChZlRiSye1bSPdf9LEswqlkugq8wgg9rKZVrCkrCsd+coU
u1Mwlsn2WoSW6aiBWi9FxlM+gbQsa7Dg9UtRRKD8y30hcEmcRcBUD4xfYut2gDJrdMOG0bbcbnZd
EtXQ9Pzg8F14q/g+jYhQcyZlnqqXWgsfEv4NVrwD6NhlAIcZNewputTOqdYwgfWUp/VTQRKvbePZ
zMX8Om2mwn0j2Hc+XyBOLIjeFMw9+N9x+PcduGyStLoxfFEib6JJAOPRq3FWnd/F5R3nA73KpEL1
PKChkXEXHOfea1q/Hha6g82LNn0OJlpt34hYSVlLCLYJQqjC/0F0BVx41exFnKaF7Qw1PfQvoM/5
r4zG+z64QJUIIsiNWXlodm5C7/kN2Xy3Sag7gaxa12WmfnbOAmxs9dNjat/KjuV9FH26C0ReTle7
Z1X51LCaXzmcMCcqUv0f/1NPodRgqWXN+bvAUkPS8G5gjVFjBdeYd5t4U7zbW2yeYFjwjIM3J8Pn
K6RaVuScrnm/EhZt3/tw378PKxFBsFfwHA0CK9r03/jJn9U4c2hoaKgDIMGXUPPvoNW67ccGP9JL
kkro4TD4xY+7Kd9f2U4m91qKdK9xAYeOQoTCCIP6GOXaDdsOy6WciWGQmZK+/rdj4Z7JIiZRijOa
vEHmxausTw6IJXvHc5dihTVOmGG3qWGrhUhYLyGvOIiZHcUBDg3/ioEcT467ghu9YR0j+GGO/sSc
1D4EIKfTswTGw+WDt1KxXMFY3uDCxzO7R6kQYpgJVDFSVanlvKsVBeLOEnJrHM4m7CsgS6TpiDdc
2pN03pEk5zGFv1A+bPLcGVX2LYSlKJzSTCC9li6KHRfRHzWOPxGN3ClX7h5H+psoVs5BwFFBTovx
1q5OVrGld+bRJWtVZUPrmUI9EJXkMmefRlBBzQSndSbeCtrBBsQdBpWyr7erp3ndEFrf0Z1heSm4
wPJgSvGs64B+0ctoUv3krKoQAdTnwmYEuYnrZTAtk7MLO7gzuot2u6aLcPE94t0qptHj5mlz31DG
4Ci5g57wyoZt0izSPQuzpFdjhNyLCfdpDFzOzE8G5p1W/XSRocY0aoF27auDE1VsDQazNoEcYYnV
NMGbeK7SPEF80YQs7+VUBTViwQmJWz8c/Exmh8Kt2UGbarlWzicDkFfUmxDk6cAMxRhSqxPpvcge
YkVb+XJdFswIPqZfI9fJavVMI/TELb5m5ybbolNfeEDNWPMn+U/uf7Gd/UqFpy+CVJXV+yGWEQ1g
22NB0nVjiAcUNG/lukb8udcB2Kix2RXhA97sDKN+oUpcI4CuKU+o7fJqLbeidAveMllR12tfi9L3
gbkLDSNo+Hb0mtue6TS1eUvnM5sRCguO0lRXTMKGJYYyIa40QSejsUClHwnakVeTHrM4LfxH3cgI
w1Bw5Ne9FpIPz2I0Z6l6eI+HZoU2xwel5/pkAUUbDM70TL4oAxIryV7xMX072I7XD40OOTaffuUM
cIhgX1a5YwqlQkvH4wGRuuDeFbLxs96Joev3MK2qXvCwuN0ls97Mf87rBXWHi/TgoxxUGqrEIo1p
JeV6BQKVMlrHnLDiRxSYdmkHWvK0LQR5CXR82QUuhUUXLDJ+ikW+vQmU0Ij39NsC8HP0/u1dCfQQ
8bQBZbCALa3hYY3TDIXxVbxwomgU1NONWMj7+l/IYgTQ6CC3fJanqOqd+cKXvEs0zantSlyLafiD
rGdd2/qwycmwlC8X6Gvjlr7iRS4JQCUbe0shoxrXa/kao2JUDfWjbNUdPaH5cQLPxXZspN7cg097
T+uLW4TdVO7hdC096rGKtpPdthNVhBpnjLPctHtreLzYqU//m1XeLjEcpWhfC14VXGLUP9gaRiZE
j1vzuf2TaAda6ELcF3He87OazJ9M6rWRhWt57IexrLxUl0UAJXcetWRfgbeYsTm2soOOeOtsJn6j
IC10r9B0X33cCwaHkUvW2E6nOFsQILPKexI7fMYz7vQuStsubilrygqcbGD294pQUDifeCEntQb0
shqTdYE3ZdGf3W8KdFVTO4JcPklPH1SAcKshYR85Dr1F0Q6Rau1tVy0jAsIGd5fN05aO/bXKQdHM
zlCF5JQ0IDBOx1+fhk61l0+FISa9kQzZOW/SeoTmX26gK4aWZ2ApN/1sZU0BPTPcWvtTdiSDZtgv
EFLZTmuEumfaixwXdnDmGurECosrtqPxj0qiRxhW/zFkm68DncEQS5fSSlbKOVZzfBhFBHd+j23M
9CSJwfsw9OhMcPA6zue363vXlADBqrhW82ZOHlxBpNYc0cQShobVslFmBb4tUwju0zJ20TRqSw8W
SuUkmpoG7i92WX+gMfYMHoIFNKTdsyC5VsyuAY/k7C/IpGzGTbuNbSLpBTvk9rC402mJcw9JODug
hTfKj1NTvSw9HdJLRzrveErb+WWk8kkScgWr1XK3JbD2EsW0pZE9IBGNjhB1vKBNJnExswa3nOlt
UH+t3CRdFqQBTQv9sFccF9NqUmYgpqUO3QifFuFcPPM/O+3Wz27snZuSQH0piNfMbmniS0rSoH88
u7aEPnzw+S7ye+6PBt1GyqIaksGxUiUOyMLEbVufWVtVkWy1kLaubCbybdY94dP+gMYi4Jv9xim+
6l0+tfO+OIP/K750PTqgIEjeCGh0XnnC341am4e3ahLnnMgfvhABuV2ocotFWZQFoQ7jij8R5h5u
yPrs1E0eomvk/TNilTj9zGBvu3J/vDbw1emItEfyvX7t7ydWtoCSnTc93VnAIINl3DB4jMQTF5vn
8+KF5hvkGl0qMaqk+fnNfNkTTN4Z30Mjw9TaF7Mz6Vi+4FEIoFyM25faEQ4Gu09nNCUFswzR479/
4kgS4QDGnngssRvrCFVG2+PLIGL+35sj249cTPfxnf+qUUfHe2VXixuF1eHCGiLyG5pSCZuNLrEn
t045GLmVQkkLGKA81Doi3n4vkavOKrBHmJhijTK6hVNYvrCwaW3KnQG6zySyE5amqWhsc4KtBllY
ZWmme8rLP/HDIso4T+MHrhiScLkJ7CZxDjQKpN6NrDWmILKscIh8TBRfkL6A9v6y6M7CGRoiv03t
2cecmPjRTFMHX7ioPjZLEHXok/imdDPgfzy6IwtJIL9wWDoW1OkpU+BhhgGAbHH87EoA4cg50BK1
Fn50IFrEhedwJ/Qw4Yu5ULa1WarlijwGmzoDRl2yHOgHTZmrXA1AroORndS1gbRCi51EWhT1nSQc
vbw6f82WQBH5vQfFJNRdNFyLb3dDB9qSleLUlGHWE+MNKIDPFlyiD9SyEQHtp5oPFuGTyP96ZDBs
W886AwPX2J02F0I5nUq12MLJfR4F5C6AreDiRwxqDoiohrDAB1OXGs92o0QqlEcyhddG1kJS7sB/
TWfnoD0IDT9rP8SxH79ZFxr1zd+wUNf5HaBZsksGKyC0Rz9DCZNVOFyEo8zUaasxAf/HQ2ce85rT
EAimoIG6NLDzgp9KnN4CpQbmvrJQQKN8JotGZxUxnUXzhzvhX+6+/fLpJUQQyDHAN9kzT2Df1pr0
Ycy27KQFJxwtHONHTYXrwaE9dsJopmeEtWNtcXYDWKUstGXwwUob//ZEmyfUXfs0DpTKVW60ULYK
xP/pOq8LdEzusgz4sorTd6QPJ60Hc7v4wqcXU12pcnaLTBccrPFscdjf2FZzrU9H6U+D4fIuOok9
GZxQXxKyA7GIR40v8K/VV+CtYuNmB98lqewZZb/9Dxgadm1TxvD3SZBpr9pQY5wpzuFRsmDP/q0B
u4/LVOIGW08cHXZAXmNp6Fj2NTR51WUb0TLIdvVtR7mL56A62bBbS2FMyjQJWA/DB/qfuzN/bMYu
bhUgzYm4GbQFBkpUbjqAvgkK84966up3ipebO7InK9GAqRrhELuzcNN2yFq8Cm6zmIkfkO3lqyVt
W/lagmluRSVbRF1xO6NZuX42KcF4ST5/l1p1X0+D/+EA/uFsRubDBsHZ7iKfRPTD/ERPCE04ryir
XObruGDaAM9t7/c18fnRatJOSXdvpwONmL2bMjJxjylCN6vUm4C1BzxUDuW4E+aXhxnCGFc3Xarg
fbkiFgJjep2iARxFLE/69e74vofOMcE7KIM1LrYrVJmvcddIDXztW2os9Kq3tT+llBn+5hG58MaO
QoKTJ+fDGSIij7SHNa3P3DoqwSqEM/LtC/AtpxVm8efTOpzCB7H/f7KZuKGvnhCMaWy9yYFZh+8/
geK1PlL/cxKhBqPnEYjh7qOXK9t8hyz0ZG4j1LtpAw1ntudN+jjn5mFbQE3PntM5Ac4ac9rnL98S
sDzm/jozl5k/TrNmP3wdJeMvVLgAbTUbzIJivt/CeRHsOOC2gArBMGsgNb9+AsMgoq69P7BAhZ3I
+7VGsXwwE1JMqQKCkzjbBsffIDRghZUgDqQb67W/bUbDrkALW3wlRtTXRFtA3W26CYJ6Aco83tF0
9P4UtGTNu7ozMpx+EFVuelA3S5GAn5LOEJO80FitafDrvD4LRGqeoS6LY0ZxwlMM+9neZ7NsCGHe
XbJhOXWD7/gL46IKt2/qQOSD12zKMR1OiJPzCQofiU96CBIESvTLBCeKs6o0+aBuwP8Dh7rIWmFJ
tuarGjEu8cNLH3d209QvC1os9CAARQHV9YrMNoe+qk7XFn6A58Piqp13nfASFZpazJHZcR0oJWl/
tLKIq3W9PXqUo07+OOxOpkoY34vW6mKlxR7JQmsOTlsguoC4s1CGOKDDbwD5TTd4wncSt1uyziR/
7gnnHZaZz4WPcosUEzNjZY551wM0xBCbeycOAKIbpZ7I+auRKv0il3IHvrr++/vbz6rVH2RkN614
IIUG1i/mDguVK6A9yxu8534xutmmKu7ktK00zHwJn8B/e8G/kIjwol1OfQgf63pfJGaSwz+ziPde
5Zuz3WuRuzLrCcy9+89ujpM4VVLWEVlNbUO6lwncfDB78AA94HOw2quBVysN/udQAdSetVbK4mHO
6V6pw56lDdLrPT0I/30xQZ9B7c6f/DYO5URCuuPAWUGxL41HtCWTiPxHh79ygpo9Idq7VzFR7Ygr
Z2xB573Rim4KxdbR+Bp3f722HkpwZSrg4ICMrk+/F/i5LWxIaGHNHTduhF427vs9JvTOmZPNVxo+
R1MwELXfVyZFWXUoiQ1K8EMI2kr2/kNKs7Fa1nzsoxDIB82yEd1/pzn/sCopN47quLCYm1sOjW2R
9UjUX5o6Fbk/88A3u+iJJXqYgd2GCk0pI24r4UgqLC9owFOkyo8o1KQROydWidIulpED/oxvRd0S
FeMqMcSLYQfkGbYsT2fmM+T6I+DExaUNBMlSkHR4rbXsq6IOZvF9K6Ka/mn+hu9vL5YEoXXKYZx3
NCU9ryYInCIpOAcXzS2fbu4VYo2zt6jqd2N5hWhLUxxNGgV/9CkBiVjYqmAvutNEQV9yQKmIVbel
JgWIrXg/VgDSGRCO8rmyCrUX0MuNZQGdN8hlCUgb/FMhtM5ugirLfCQ8C2kJ+/7j/Hb1Rjtv7c26
K+QoyiaCU+E9veZXCPJRhRyiqfv0V1VWMqzOU0mZUTkJUjo2NlyEkghrpP+P/ZwbqGttYC+22heT
nkE5vGAnIyoRyFsyxxLYcSFzOlddSVJaw0596yd5sN3aG9HX2p9WpCzlrdtQtI+umtxN3s8HLKwT
e7HjUUGEQs+QSWzpOaglJQXgMjgX5tJbpmr5EPfRu6yjJ0f83eLDtsAx7TPlqj9F1W1RIwZxoot+
19y7koEaxIwZctKbeKKb3vXIaeNbulOc0ntzODqm5BPIVC2Z1yR8frU3zZ6n1OGDj/0+BxeCYMrv
5okAW0R4e0WH8J8Q7/FGa2eA11yJdUkS5t6GWvbybRsSbfpIgERNOYz9C2RUQwsy20N3vXo8Uysd
CaKurOwuuHeOz3E1ACbQRMSFzS1QD1EPkBAxX1HOl3Q8ZNELFLjYQrgY4LdO5LYOnkqEuMrmJMgv
PMhB/wzXApo8hKRM8U8Bm3g6bZFMW5oEQdIXWl4ZlHapoxnHArUn178XrDlier4hVzHPxXO5cQn8
aY4mOa1U7XYzAVX8ZWVnmoVfaiLi37S+j5bTWbM7Ry3lQouvbK/V/+SNyp9to70DA47avUFxoRas
8rraGJmKKcvem50Pcdb8XqSJBktilBKpyEgdZVJSXfRlRw5TyR2mJo1B8zBH+F6qpT0htN/9ntzq
iuUgzEeziMfdqQngf+2SH5yX3eCS0ATLC1a9xhu15u3byKaJQ+g1izS/s/5gRtX3IFHPi5AyMv+N
i5FuUuG1DWhmPRvrxr4JL7O1/dLM8cPtk5Nl0Wy+RijoPvzFRIXFqLyzZG5hACMes0tNOTFWrP2i
p7R8w29Ylw+am5I+0hW1EUwievv8HcYNeTiSzMKWEn1drQWsS8hARLZI+wuZgPkzHBe75766sC4Q
MguWlhz8iWL8afsEERehHNH6JcO6OMjLGorWmWHHeeCcD9KqoW/vJ5I7kvbUsBdPkxInPjfZNWGp
H5w45ywsWI9ZnMj4Y7mucn35USRP2+Ve6LzRTOOa44Hrj9A2AkZ5+JdqoX5twBejzRAUVHw1imjk
eg2EuNRDjJhBSHVOEuLCWSpST6qAsidk+7LoKLFV0qFOffKt1LBAnlRuxRw1Siy6ijJ4xqzG1ha8
NE70sQTP6MaAhEGZmffE6vGYJwKkRXqQD2JabaeZTSY3p1vD0KT8QXrmWYoNO1Y2JUPoVqqSbYrY
1nzYSGsM6e2rOKQucnvtZX255LLlyeYCT3B6yg/II+JtDzzrkz/h5zSCQqwyjZ6JZ8I+58Qo4JA6
2F6pgGAfWJL+kk5pyOfHO6pHMrfGe2kMAohsLA+tU8bQmB9NyjPyrDFt9IDYywqCb4bxgoQbWMry
ibwvBZEr9KtWpvkWdpHlQ3DUY9hZi86yCrKHgjeqFF/VbWZ+QrgtbfQBkOB44bPuFkqTURmNfXFd
U47ODpi8pSoOlwgAuizV1oNbTQA5p51JtF7pFmkSAG7bF0zUa8VCXuHLloFMhPl2/kJ8WkD8hD8g
I3JL/wt7zamtRIeKlsaLYgPhDFbQdP+OCVJWw/7SX8N5hDOvqgt+SFM4f6ph4P0UWMXSJE6ObsnI
rxTnTUQZTHK/KOZgGGXelyCXsE6UCv4J3MYJUNGh+EyQ3V5pz7vxOmpFRLUZjRy4/VjR+nIGKHDM
1/Al0HiKLz3HeAiNZ2pLDW2egmxsOhjuvkpJojJGZwYVQqU1RWpX0BV/Mn4tyg+GV7JihHxClXwW
p8+GkDksfkT8ESjQjxCfvjFB3gpPDo3oq8OeuDkuDxQ3J1fPSyjXIbeb/4znbqj06m5VN/4Kxjc0
SribzowcyDKSbLQn1EkIorVy3VEkdC8wcc76DVLMLx1TwRudIUgqe6u7HT2mdSmrQT/vHfuzt2p/
BXm7R/vI7ry29UJdeIrGxb0zdeS9nKbaozmYRif0iSr8ehf1jeaMmzBD51lTEK9P61drsbTPviyA
d2X8D6UOtWm22G1/2mPpZtciUZUWr1bwhrAzw81KDEQJiQtXq5bdHKDTi+PQMLz0SElHwz6VlKva
kOt0cYFSSDwKZz9iEXxTFclq23YRymYchbZyAfYrNdUlTUy+UP/nveRmrZZco2refMQHYWnTSkzX
/md358y6HBEsKaJTMPmU+/EPeuxziD9u6ILCDy11Os7huXvWwRbpoMSEJv4IHRK+Gpef6nUX5AQA
RWOQ8VVVaauOZ7icj7eQJCAEIRtR5wGcz5smUl6cs8R9Kx9eTHDsOuFnEUfXLPJPcYk2olR11DDQ
wjbI38AG3lsuW5Pn/xUOGf2fMVaeyo3TN8eTtTo6fcMzgBmOUNa2tVxCes7Do9qPTlGj//Ed5qC3
JATkwL3MpYD6ZW5mhCYCChDdubAEE60pqh3F4YeFGFs2tO4SDWTy9eTYz3bx8ffAkJuwiOA7RH7P
AO9gRzmsrPR0Tle3//E8DRxxz8c+qq8gB0+gvmWNxCjpgWCUq2UbJPiEz9vHH0ZwZLCOjfu0MtW2
2FYzQp14MyUL1Fk1tnwjSrsZvgNJi3S2uHcVhBuVz63x8+LumvLOlkH/Niftbu4LqwC8I1LC3Ur9
n59VkNkE7HHkACHew1QPYKDC8RqeJE4aj6SpztXymrAtFEHXMt/wLEfY+eGYhJj97RuCwhM0ytmE
j4Qs9x06ea5t5LV1mENuXkp1yqAY5yk4W/cPKt/9auz9VnL9gXbgpMZH9QyYQrUaIBEXNuSH4o9N
E2v4veNmbnwIBEeKRqXpdwVY+bgP+g+neapb9uZk2uboqFdQG81rOLNnZFmhlYqogK/Ot+2oDQ5u
Uqi/do7jG6pykLjmBc1bL0kaf4gcMqxEXp43LFZarEePOJTtmV2D9nG+XGJL554+oEjjeWcPG9+8
NIrWJB2n0BY29jGR0dd+IVGyH3MwIEuLEUwzgJmtuaLjXMqYALSf4Lkbu/pnH7N4l3/AeLcECDOk
B3YfITnAOKJ7ZjYUWoTjl4P9hAvJ9482KvnrRZnNaedOzi2oTa4X+XihrGYH/E0WCPFImhQKZC4Q
qg/yZrF0waaZDOHLjqSdkL4/cNgBv6V/tMuz/EHNNCWcDWd+k70IjHG6Dbfp99NRD/T/4H2xRFtJ
Uqi2Xkp+HaIFgPPp/MoQ1rqVSeXfuprjLblMrn0L64ipjN/0/6B528s3dOlTOob+tKfUsAqXO/vp
oTkmomxgx57+KAyB+6fB9m8M/8ElrqsIL6QHA2nkM+FtBirx84XoTC2caIDAvl2cLPBIEElwvzTW
/TRpkD/B87idh+m7U5lTbJkRsWJ7sDTBAEgoabfR972FjjQSq/ORaI7uwHtAuCwTFKiQwgJHjxKj
zZip6WrySFsymDp7xvvAiZdi92mlD8y5uVjL9ekVgGWezKYQZAO64EEjs1EQnmg1ON4mRCmBJ//I
XV810WtmcsWJn6DPC3ww+sha62Y1EKwnP4ULyLUPcGrRrfgF/uhYkjwOFKIObr0uj0POjkoeOdA5
9jhL/9K7vzXFBKVxIEwhW2gA9YLpGR6xWzi90uv3AgHMbP7+P/NK/Y7GhX4PW5kHivdjyxAzE1wh
+fMKl9V8uPxDn5342U88bBMoZ4BbetPiPl+4eXbroXbAS+qInbd+bCP0zoKyjbBC3ZiJ7OZgpCsw
I/xra6WLvuWLIJULO2/TDDaPr2i14Z4XtF5GQxO02UN60MS0eKYeQt8gUcLmOEQuAvwkKb+groyZ
T7ZXBZjn/PEJhNMy0/LiNbnof9OYs4qarQyg2cZDfm2Di/zFKzkvlBZWdej59ahkkLtjrLWB5J2m
YHqNMrESO8W7iWR1WJafPOoY9rIEl0pQEto69d90U1+vdR/3NpjvtBMluCbl7c+/Fref9qd7XcyO
toj2g6R2w+GrjqifQ3uKmzrl5V3c16dtzRxvgS9ZuUmDO9l9CuKwAObwlrLSJAWYkCBq26ASQX0A
C1C9fQqdSOuZDR3WwRAeWqkRoAkUSousY7D18yTAkMjULc5Gm6r0FbWFJnIPtJh1n/869iyl+qyX
x0q32DxM1e2kRmZNQ3iiGhVzoz86vxsFpWTprat9YKphDITBq8fjqbRjfFqksFAuVAjXy1t8eqj5
HwOrhgIbus7FrD/DuqFMKZEbG9z9I8BL5AMqB4j/MCfe06PMzoe9dFiwAkl0+9iNB+cDhW3FBS3t
EsOZGRunEfwglwh1n0Ez+LCj32sGJ7hfXNShS/n0s4RiPgjzOaS6JOWyTlvIhQvdHrgSlKBiAhX/
x4PPb07aMQpAbYt6f7lq/iZW4ozfk3hTisT3dUBu1Dq7gmS/9rNnm76j+XwAJwijbSrH+MHI29aC
rC23Zp4Ymc+G3RbxXPDwpnOIC4wsxKq4JIg2ZGvZ18Q/+NYBpQGt+ls5kdNh1nI/MQ86BXb7m4Qy
gM4OyuWOC7vAHRaUcz3XSRj5WDVpCqiU/66pOj1yLqNgtQbpkueG81JkLabSNacdV/pNNhvQZWm3
s100oLX8loAgSn3FrOKyEP3+KLXNMV4Hy3NnOrJlHEKHytyGu7utKF/Ncq+/+3aI0HzhCmAfoItP
6utZjZxcdCD9LdVPytQ9QvMT0tcK2SEwF6zjmcwusP1c4U6sNAYsMVXZpNgFwVfc4YWKe75QRvsF
864fBWn05h3aR7E+4xQfTPr2bgBZ1A3nxaEk97sY7V9x+WE/i0xByvpaLUq7vt66/YmFahwv3x+n
R9VGPGPxySDE5YvUuyvzTVr8gAo6BMH0la73zzGcxFv3AD9x2YRwj3o1J8U9B+dxLt9sEr2RN47f
KJPRE9iVdWyUHQBE/vuwZHqNjugNApqp83MqS1pyWuuVXkLr5GwTUcachzxlpOnWN6LXkvm88IPk
tgAV0Eodb8r1AFSI4Un3nVHoWP2vdciaHg6hGRtgjvCcZO2+KObetMy0bfld5l5//sA+Yo0segRm
8Hm/Yqh6QP9TOZ7QGGysxsGzmv4RIgHVP2ZVsmeUQw+HdlDByTxM01FYgDmp23PUvle78zrX2bEm
nGV0zS8PnAlIWjf9thJbyJXTIZshz8Gfx35QWfMe0oE7E9wGJyuS8O8/7xxnW5xEK2JclnuEwgVX
P1Uprob7cu/yF6sCfhKQRk40Bg4tpRGvgGYNK+tAYGB/z+fnMg1qv50Ee/i8B8up892UqGWCFM5q
SctG2HhjdMgfASBYGzkkkb9MEBihuBAbP3zLn7PMHTqRPlKyC32tt37N/y01g/XZUZ3VJwQF2czA
yt+j3CdUhzms2eMIL8xu3yRS2nt48Dc7VeYmvZ5qXGIBS8YA1BqdraIl3Nrb951+kUbZxVBd/34U
ncvsIiLhQK8T/0kDRG5E4NqiS1Ng20QSPlDGIcc5ayrZ0i7jbVDOvrZL9AC//hDivnkCS3KTu1Ff
ZwcMd5uGfkYiKh4Of+scb6xEIigzZFjNXY/K+8Seb4SZoyx3Sodupw3pQVewK1G4rNptq9gYebvR
x8ybbCtM/kumJ6hF3MeXubTpBqyZSwRgGCI0vfHzoL+a/9zHZY/DBqEv5Z8IbqVNypGRp8obQkcp
4EN6pvRD3rKT7pq4ptBxUa8jDIFwW5Rtq/UsRjnpDQs4reC/dfsi1OLchys381Gl9811Pr1IbSA8
QFAD8pmACujeZrvFRG5nRSZmXPtauBRFzXN+mvuAmRUlhok47IDB2mTLlTWf9Q55Zztpr82+ifej
NiHFUd1hod0MvMz6hitJ1L8lgSVp1LSRCtu+mgTfuY1BZ359996GnBs5Boy8lyMLuVWG5cn7rggg
832GuvUZPgEFwRF+S/tMeCeASZkCGGuokG2MAWUQM0sgp59l7ra0PymRYUYXyvbruQICIR1+pGWx
9FdsmEaQ0rQhIFcL2Ym4fVQzRu2H1DFdn3W7U9ysThZe1ptQMFCgD9mDYkPrK/RmnqII29attmO1
3LYDxnMnPo0DmWK20dqQedxjeXwEXvqL4WcFFvE1QR5CrT/FQgDIv5ZJfnoDTU9mYX/VpF4TdScA
vRPDU0SeQ0mHLZAz5VN4r3aOTfGzs0DAMuQqQpE2S5LF7tq3yddWg3BpDTFV2z8C1Yb9xWdaeeoe
fajr/hDMiJpT+ejq4pqskdgNOziLiUd3D3BcBcjrkRi31bp/MusrbClCsbtZ+ztbK0YYF++eJY8r
CAP+7qhPhwfRlWlKe11ajUPqdyMR61B2Lmxl1uFJqMiBB/vXDgBC6QusC8G8o4GSWMP9qV6IuF/A
+D6+yWzQJjFozeJzULddf7VzV2CUXwGiyJO9P6d4C8AR6J7M0WUuU4kmX1ZgpZwTg++uUpxDlhdG
SQn4C+jCSlbWmXi/D5wgWf91y7nTN7BEqeBENty2TOSXTvsTTMVi+cCmua+7IVREQO6dgvc41P0K
LRSWt/fLD4IywNdUc7ffb//lOasoCJaZuQ6oaFzcMgmaFHbPZ5GX3Y7fUeZy6O0Z9rH2uKUAFY5i
3SCywz16KatTpglIUf+PBDZCaPjpEmeFgsnQbjhtmphu3G05suavHlgQzauG4G5WM5RzFavXHC90
pd7XdlwJa+XPMt2WpxeDByt1Q+eOQS2PS4Z+JOTukfvIh/+QooQJJJQH7Gq2Jp4s3xP9OKh8KPeL
5V64j+ngPk83K+SXIoQ16Ff1t/Fr+turzz2kWL0IvHHHRWl1QXXEI8tC6J7Md7Q2DYF/irFJU7FQ
NkInAXXSZsc8L6Jk1YSDV8pziKDSOe2OavfXkWOWuErvpWnOGNBS9HqliQZlUaCYHC4/YmQWPsJd
gLcp5xHLp9W5RYSrzQS/sijX2kbKlk44y4VfNBRp2+4f9CD1LTNlgtCVU7kapTKDDM/UwYSu/h9P
5Ekhr0y5Z0RkOZJ4G8J5981wwZqVvhxJXpaRYC7MV3zOCpkdg/JlU78q9XmlVfihVYAQbGl777Gs
i01Lzj8InVCpg/CuV3QwNp9ZtoGShSuYJoeXcp8KTbQSSl0KRG+V2ZYVQ+EHPxypV3s6IKRcvBHD
KiZx6/ESoA3vVHiNKrTaZzwnJBYdT2fZ7ThzJb4mmus+sTOqXzAWkFJefujq9urp/zLOLif0uV5J
rlE8jSMdMJRlPz/e0XQeL7CCzqmNwAS0/NMt5Kvz/27RX4XFPMeeHZVRYlxmxwYxPynD5+E66wXl
HGlaSyJRhBaBQ4UzE/ATLoQ3sIxh5dYOXjFnVFZYdYDr4HHOyBAhwHZeb4upIl3USm0qQCyzZUU0
W+gky1T0S6G0E9zAy9Jjnc/DcGz/evFh50UsJTVpJOzKYW51nYDEHMKs232HVo+v0eIoL0cvDYK/
pbd0tdsRNPheGgzV1ZLRqqbK9zxekqaE/+C+XfMxNCZq2qGIPuUAPNPyHfEHF8iFPHVPigCdfgbE
8mWR20xvkZCaucAKOKSX5/QKOEabAMeE8xcUepZxQqWFfyqOCGqF9ki8MXqbQP2osy6TTWJi/cEE
3hzXk8infJ5oGbAINuURa/Z690MGrFi13XL0LUDJ5Mm9dw5lxNMRAIxKJtigANmfZ9R1vMlU7aUs
V8SiiNyBlStzEXTTJXaQ+1z3w87ndEUfEhEEjQguGLP05iNIGiKET4QqyVBx+kGYw6zWe2dtta1y
ivBctwjBlYHX1dErun7tSB/garK52sVxTvFSZZ1F2JV7RXnbi3LLr3IzNtR/opIUa+b53eFjgc+E
JSppPvZPsqW0MZzmMPM/mEvd5P1D74/pcL1r6Pm7BYfFc54pCQJJE76F15fcJkK1JYFQddZ+CTI2
oPVMevIu8fzOdLIy+PNE6yeSel4QW3acxlljn4uzfD2wb//9126jToIzx3OGWObC9x2lL2SlnWCX
LicgbtXVlhCq8reGuX1RrWShkjut8Uqpo+SGLqUU3xOnPGCaMYJi03X6x3KyMkf+upzHS+MlUhfU
JjwDdSA71fObHGD02VuXX1nM09S151TW3dPpBwi+5YWVIdnxMfLQDoaym5WKpR2rRwhAQA8rLz3T
+pFY2jSlAucunzz8s3nfV5BtT7qsRzBIgEb3K/uCv1OnEdgqJX5ocBcCDj3/l3ZRZuBjxgTi2vW6
ZzOpnZAQWRKHGZA5D8gUJRK4Xv7PTIXnE9dYXm62HJJnaw/N4aBQEYxIHux9qzmE1P5SiUuoedzi
d5Y24Dky5a6j51qjeDb6Ur4tKD+HjrxcMPpAg9yoagEOgA8uKgaze0UlGgE0gfs5Hs35zmU68Wwk
vjRGU77FiR4pOrvjaf6SsmsTAiv4KNIeTfd+O/yaOThwRMtyqjyuNgGqYFNeUgLwxvrhlgWiPeHt
7BZTu+YvZE+099zV7deXsOzAd0GQXw0PeLzJcWAZ1KcL8Cp+/dybAFpwqJZouv81PFhDMGWt3j0w
DbHl3L6V2VMjhRSr53KwEnNcHJBlb8BnZslGlLpVEB9QMozkkH9lM1hdiJHvjwkVimJuzz6sQv3N
wKTkB8gMvmoq9nqDMCFJfsljCn/L31RXEyw6RrCvw9O7XoY7IZ12SrENycixJRrZD7oLQX/V/mDb
WK1Ir6A3xzA4fG8QJL9jmGA90k9tdKtl0Mri9CsmCWlqiUjRQqruggsHpqQbFtWqaM/otY4olGdX
TVFuphyoXYA0yRTeofDVS+kwdT2xMbM+wpYk3E3CYo3BFps9oZdjMyeWiv2GPW31FMqt8IqWOlvu
8VvYZ75GtjiSF9dfqaMjZvZCPS9wkVVEHLlpycMlv7yF8JjTbdnMB2zL1YlefOR4ir12syfj8QUB
s6kottafcb2dkSlvjAcbAuBVdOJ3rQuZxSjwUulu5z3hClF6EGHS5bwI3SncB7+dtHGcTlhad5jN
/6DYJXfwD+Y0SilC1b+JzzYWhbRDWnJzLs6GbVDcgJfw2CsDcn7r72lxXpuOKckpJcqOVcFzO72l
SBcq4GY2QUaPqJd42KqE0OHrHzgtByeyLd35zTxM7oF/v7mPhOx6TDrm6OZjbkCrXr4MOmaFwcQU
dqRbh1AIvUE+78hf/c2ldZ6S5WwE06CK2bdS4Nlu3hVBtgXeHCgyjPZYfpjvbJNBV0ID4E+AhjET
hx+v0erpYkGJwdyUyDFkBlCdqGebq++h5DoKe6ZEu+PImbTL/h+jXXR45XLnurQv6XZDMFmaUTby
R0w/xL+WJZGxqaG+3KEFRt6DmGI4v50yyGaQEsXzZT/O5Nhkv1gehTZUxrmnY11CIIHPQPJvfqHi
XTpI3wtpbUhPM+rrDk9lvysJW4E5OlkTsMoREq+2DYPJuaQOZms9hqzEU4p9/HN0TZcDhsbIFO4D
fFTvd1wPcdcxsS/EAhbCXuAaG78LBxuB7fjK5YD1QoT+1+qQxUhidydLHCbDntV1pqt100JAFzym
z+9ukEw7fZeE5AG/D8byXlKOdyRzhje9aZp1+AxTVppA34ppZ+adrhc7Rb77OHVLGUWmDYeObvSB
ZxX1XtkItLvtBD/kQgf896ENYOMmci+LQRLbelzAAi5iuveo00HuFMcbYa9f1b1f1sxYEIc5KPkZ
g13+Fib0X+OIX+9Fj1eXJTZPtxX1e9MWfBR3yUtwVyboG/wbEEG0HNvmJqBfmJtZTQTJJNR415jK
3OaXeCDlEodZ7wqyZBOFkaePDpdmbN7DPGVhtdKoXN1U28o6rlIFePuHtNUMaKbHhen9dJ5itB3K
YGdEAg3SVnwFLZjyWHjd8SSZf567LJjYQcP+677ScfBmhZcXL7gCoc8hbrw/lBJiF6wBayxTOTHM
WdeYKerKmNNa84/wV4/Icy3Fz1q4fhAGS10jxQxVj6YT0oRzfgSJlH3TwBPBz6hd4hHsqoqS9UOW
tto7PkMPeRF5a5h5iiKU86aq/FLg0AnewwINxg4WtLCW+Uall9+W/ug6yOUrZT+1JmJImk9VpIzQ
JVCLQp8L3SBlxEaP6plvy9z34uw+k6S0pQ0CBk84oQuKtbumySwYmkOsxYPeTsHA4IfhEY0u9O4v
Tb/NWKddE4+pm31lUmhmc9scn70lYUEdLf2jKk5Dh+AZwvW6xmRF2uJiH3e7w/6UZaaZgv+e05Wu
+MRCriEVumGLSisGez3F1CdsKhwTbijVSqR189vSDqGkRhNCzDmPnmmIIfW0P/5xhxd5Vb9spuuJ
ExFmQtvIc0x3FOnzu5N7BUeFh8OZoTbBufD8ukdxOD5pzO50LiTcjs1y9shAspf3No4O2e/cWt/i
Siqqzvj2NsovQNqNFdTVprRbzl8WLuTL8BBq1KpJb69ox7I7imVE461MsdEVyGPPNIhtGTspA89d
NLDl6Q7A/B12sJnVwQbF6Uq5LqhApru9CQrOdbg1zUeDZ6PuJ2ZAGdRkGraQ9nBovGXfiHT8q8Vu
nACdedzPW8b2Ulx+UTmltrJ262882ndDeHC2fqCNyhaMrVKQA0jLYPxtfMfER02bgSs6az3SuGHW
9W6eUeZP8/WQe2JjgVKUWcqTQLCMJ9DOvhvFGEdN6S0gNqSph6btFsdrPUEZqlgnqpdcqxV/bDF2
o9pF6pyuswFuZZ2j76KrOnQx0inmvqWZtWCiqAxsjXpln4IK0YMDFRACh6ELMAbblIk+m1oZCLuI
lg5YVlvEBSTxmYQ2nos3TuWy4chZSRenm1KYC7NaSlwszbD5BjRRmpNqd1lLbCaXEWfuJ0TJIEdN
H10GJJat5McacU6LCw3//dXHoA0MNZaS0nhDOEIQSDDBXr/Q9o3fcNlcdC0ux9TfZLRk0a8uDT6f
6AipuQCAcLzaZLnxZzofP1ctt24odlTufMTVtDthcs/v1Fd0sMX6R1HAAqIwUJ5plAAaDKlXOsU9
IIJ4CuyuUmghCRWgkkZwwcWt53og9IDKrbiFOVsQ7Txth5ooxecehMR+X5eea3tmxOHmjWFhXTkA
0hIy++W8p3SRlbIbQC4zqOdWFnLYGKYnwaGw7l+rB5du+guhfUD+ptnZF0jYBKvQvi+SCtiosy0L
AlCj0jlOA4EHVRdjnB+YvL5LhnOS74y0VaQBJvSJufoEYjnHONHo20D6Jo+HcZJY4gt8vgkMq11M
UFt7zLtPT5xnD1DmtHrtfSs/MGRb8pfWNqdCgIhhWD4d2AtP5CLnfL1RmL451t9aTguqz/7hedgX
SYtgWSFuS3NYe76uG42Cy3KN3xfaNUORYg9Ew+eXiBvltcmm8iw7zV+644ZyWEmUMJ2/T+oocY13
MeKCkFrYXp2lpBiN4+J+OcDdvRM4w2OrxQbQLv7jhexFqPXvxBLEBTifgzGBES9k4wv79H2h1Yz5
FY5aNmZsX08Ms0I119xB3n13YtKG3I9Q+GWCxAJBgS2i6FLObJxxurhLHwu2BzjBmY4ADF1ylSEh
xv/cFMRtIX4dewCsu33q3NXPwXT+OezVILkhDcrva0wrrWJeRalaYvhq+hJnHX4DCikNfWbakTmp
X/0hy1B9G2DMqtk5LtSGsQLcMCD/S8SwY8PqhTECpLNY4IMpi/7ty3/noI6utfnfPWAFOF19BfXn
IAMpxDtiMtSvxyhYxhGKR6g59mIgBnI15XMYigx6uwB7nxoPrbubVsIXauUiBtEo6am6NwyJDI/G
yPoN7+Y3W/OJGuIPeo4wVEi1cO7Vz2mrz6pkvqAeN5vKsk9hUo2Dj73w3CXeDoUku19Pd8FbWPZX
Tj4Veoa8D7ko+j/5xugnxB+0QtDN9nPgqb4pParfl0RCgYHZKl3ulmxhGCGmtjvtZ0mo1N1CTydD
ddFuENPEVYVYNYM8il6CYHpEKSF22xqptjxtphpEsPuu4rNnWSWB/Tw8ocYZRTATU8k8I2CDTWr5
iCZmDQuNctWp64bC0H0fWOqzE6LWv3v+S8ZQVYClyw1ZpEsJkt4lxfhSLupUJe09CjCMZzEO2qCu
0wLLkDMfh+yx0AdN6CgU3Hmaom0s2u0wLXnASSH3OiDbQwI7rp5AbqSKwVBwXpyH7NGliFavyHlV
YNQQk/eqDNbnE0FqS7wjrebxG5hWit2/043ipQLhjzaAdoj4aR3VxsYxNOHo0qOXqyS7hAf/wc/h
ajGT3rrxUCBEP90ghDc6fI0qgjmeWaKFzYt42fmXeWuR2mCLBVVSxar6w9BGITeGdcftfgR90MvE
vGWPtsgvREGh5qgoyo+N+A/6N3tQwCZzW4en1ZsR0d34hamSlFDsnlpMxv7wmX0We5YJMqN975N9
Nh0vEDtr1YzeJujqaDaafHEmlKiPiOUgkLG4tdYcCusL0nk43S9mLLHNw12a6VkcFEltLpRXp+Of
Yo6I8eXw5L/va+baqFjGzY/wqBDl2/ponCGAOVdSuJrxsQ5nyrrSsygeIHWiI9Nxy/ReKwUhZaT9
piJ/htedzV4+lc6ZiKs7OAOUMTCyrRTZuyrzywQlnd5HIzaaOuJ9twPI16Qv01hE6xh5ga6tiBlN
FQtqHtvb0E/S19CUN4SLautecxveneEzueRle+q1r8HB3r4x1P1A7y354ACAmVq0NAbaibKnLvPr
JV9I2Sx0OhQrkXnu2L+Pd1cyJvJNoql4StkrZRlFjE4OK/8aoWPa20pzkO6Ca83dYjWf5R+6cdAj
j64nWRGoAHMtt6oxRL/mDy76+L6+CSO0V/kyeLH6B6Rn+O6vkjix53xZ0q+4vndDanv4L43t64RR
KMcTNj9/ExxVkAJpyIaXGKLglTxuCjG8Icl//UF+SmDNTffLphFujmarUHFIHU46kIEeN0Mjw3NM
M1fHmrW77UclkaLwRwxSThZ37LWNeSbpduNbi515MnGio6XsAMGsbI6UUaI3A5RJ5PMmHZooWcln
rjj7Q3GKtSzIjiPuHeIZ+KdyfWE7UEGKtjoDJuwcjMB/U/85K+hGX408EViqVxJhvL4GNnlYeFzp
71g4YQRU2ZlimvwEHxLNRhLwqQ0JHleDzKKiBO6l2RWxqvl+y3OzKiSYb7JBPVtp0CgvaM8AR3wX
Lgcx72VamQxoFfYAvFJ/Jr6KspmFNADvcBGeHTXpEzJXg4g1i5DvBHbvhoqg+h6Yb9MpYreUq5Gv
hsNbaxS0rlVeNApE2z4Y39SYaZv7q8ukYQLg5oOxw7HxhFDlMJcVrOp5bkIMLiMcKOmY+HiCiYN6
f5YBuXVkOpORayAm+qvW3qiX8EMC1gL9CDydUtMSBWhB/U2F94f8j/fIKzE2OfpeuaXhEIjVciEG
asdO5KBUpr11rhcSBLKP13Q8sllXRkMoNF1kwH15jUnBXtZjJ4+Z9QyY0/7Wj8mNLFxmmeVbDr7B
Ieq0JviLyHjoq9imoS80fG9e/HUNX9FKNR57MwYqWxpfem8erH0mo3WGMoRjbNmso7wn/MOWDt/0
Qh8iEQ6Jd/B73e1YmfWLVkCeoaskJ8o3jZlDSBB1NG9XKdb/UDcKj+hF/jKactb924iGtH0h0Vrx
kh6R7Ill6mNodMRIIaZPzfA7xeuSWGh3uAToL15fzEzO4mtIYTe+06POn9qbcljspWqombQJO9Wy
Gbbo2HDMWmJbwfP/8les48EzepNBu47QHj2O590LV4AOn563evWgRQvTytrVqymE+CHmOmIP39dG
0zSPTXgBXnOhJVjGteVp+2zodLfeMXTKGfSTRAuh9Xy8EHHMXiICSZDHSWyqAaLSiwvRnmUJ6hNe
op/Ii+WpiDFopgXvie90iOwQDD1g68W1Fi+2NK0a8bR2AizEsYUkPe2km5IuJ5pVbUl9RPVJTyAO
vpWJojCwkmzvsVqt3REAUb/nvQTJBA/iHcwXaKMmYIiJQUznPKsgPsFJ8pd6xF05QzfGf+8ccNnU
IyuNtEDl+NZCwLKvQesteUhjFW/dFByWpraV3r3Qkl4UYMAAQBEMWvl9qaGZIIkpLrpKyb/6u/5E
RKoG26VYoDRgpaIKa19Nl3ztqrJcoOvBotwYhQKrVcl2/f6jPDMl1jprGQCtr+2x4IZ6HZaxOFMS
C3Gb3/sLAGZ8QYJMQ8CXwdjiLuF6q2rJuZ6x2xfMUD/9F5s7hJBU9SgnBPVK6s13eAN2gyefsJLK
LTTW5nj1x75h8+Ry1CVe4qdV/Ng7cCVAe/zQlQ5rjqyCdt+QhWUPU1WN+z5h005tabqtDkDEXBGM
SWcEjHGxupHubkAdee0YC8ELnCn1TLVvefSP3OFhFr9AEOQcSKQ6bKsn/KtV0OpyAJ/V48URwDSD
WA6PgXzkLxd26HHAxNldkpui6rf0Z2cV2mCRi7sWJapK2/NhGVH0lEqfTpzjKVHGzGmTxs3SPmDA
yxgKThxTuDakhSczQ2qgbfC2+AQlwGzEz4txetnqtYF1LpjkrLfasCpiGJ3hddYPIqZqlGav+Gty
ex79sddnQ8upwN2sEw0s2rSalPXCsjSH1x1uqcQBbRuMDlDShF4WJU+qOxGvxLFiI9td47455rIY
GY1da6SH3KPDZhEtyXrThJlRMOPSSaPe2do5tGAzsCMmAw7BqrzYCNmKeROs7gtb1UxBK0aWhJJR
kq4U4FeCsDNyxVQ4cIFwx4DVCRbONr3GTOyxVl5+ZLqPE4+now0I1vYFTpzGLEZkOeD6xuJFBLbo
DGI0t8vW3PrC4d+hXJexuA2Rr8QUHzi+gm8MqV9JQdYikwqxnJ729ZIoY8Kc3tZd8jz4dAEDB1JB
uN0o2C/cLCcGPr+ZDjCQunfdnSiaLzx+X9+XEICYOTmQi3kzs4LxicSUZxZZMJNStaEA173GUktC
Ov4yX168W2lAfN58CtASpG7zgiy+KWr/1KBwiWdmZJg4KhlpMf4F/Bue7ww4InlBH2LL+LCPd98u
4VkBTTL58DIlp+WeOsA/92WM1oCIzocHwK0+v+AUFhi0AVdgr4OvPY21m7K0kn0T10FADR0gT9h8
XyrCPqT/3k8tTtbPbXekaHkD5AzJ1chSxO4AXJL/pR9FYX7/+pb4UTZcDccGoxee7dWshuR0ltEr
kiy1oTcVgSEe1duSjhopvSquOsbs//mpeys6rJnEQrAPcFJBmzplZ5fdbusw1fQn3Dzjbx8BbTfa
RzcL9f7JHmmuLdKKDbEtQnk5Mf8g6xsZEiqT9WnHmA7iXa+79dJKZrO2KkUExaERkP14wmsKXwk0
5bULQwZpOHx6Y2hTjmBhIoPL3M2Wr1R6083eT9qtC/6DnWjUqMgv1ESL7CE1Ft0unOGwVMkJ6a7o
TPq4qKvnwBxcHTV6dvu1T8bcwlEq1MZjjGdEMDnGWOVx9wbYgsb5uqpEcqjbxjrgyw/vHyc954i2
U4ZZX2axNP5+vzluaAHh/MseB0hCGP1DCqYXMSc5eCKM1yZnh6ufbHIh+7Xe/ZdJM0mnaL+DGkPP
3FXUQwPR3cHyh4M9yHatV891NRMCbImrdCgUqDWPXApSnYSmfdK1nTWboB8GXl0SApnDJDDgUQnS
iPIEFqnr/D44aLGUL7I69OQSn8gEuAFiQ4q7mJjsUzf9yiTOVoxudWKAtFPI1KceddlH1lNDC6OQ
UOTOLc1xhbnaLKoSh9fgsJYiTMdunUKWF1gyBa4ZHgurTJ+Qou+Vj46oISCl0KUGfV0jQENvtjeB
NYAsvucP39DqSuHc+XyqQQc4RrcjW53LWSl98HHcbOMdLtAaDTla1nBbRgYrQJRvTZgzHwPQ+mN4
nPBo9UwFkp5U5O3wUElIPV3bEOh2UJfXrugHojo5HqvduNW/8ClJOLzw4BfnDL9iSX2Nqekd8POZ
hsI+J2pSuc8O23Jq5vuGVQnp3XzglspjOO2mrN/wNMwzGuxo+30xfHKk1b1FIvc42TKGbLP5wH+v
b1V6bLFNfhrUv30fwtR5/3Hij2eNRtx3m81C3ErnuQzOsfeNLcdAlictbWAs/+Ehsz1nJ4/P/3I2
Gi1y2m1dYDmlJc7f2zp28CLtjCY913uVxKt1giAkXCEpZ+dnIKCZ4z1SQBB84wU3YV2i3x26GjV3
VP4Ds33YELDw5GbuXWKQgGW0Q8tzY7q6EUJcNObsYMMvjQn5VhGRrBBFr1HxrFTDnTsk39IeNOrF
n/PzO65DUmeJowmYAZjM/L5ZWCtFxA0mBu90tnUtYMX2STSpNH+m97+WTDzFZG5o0j5puEEsXDFl
8ONExkxyM9b0acF3RUlVYLk/pIONh0abnVRzAuSemB6jYqAwfVjMv7EIX5hC4TWYDICBUSWAQJS+
+EM40beryYSFGpQ0HGMLIAi012syV2OPzxlJAVLe3XZE1JGNvveQuKK209MWir/Ov7xi6ldAJO87
l4n8+SsFDcRBO2ZUPYoY2OrseGXiStkhbQ3eWnuvzVsrQq8Lx78nLhqi51AgHtoPBdviXtCI7pZ7
WhLxJ6LjXLhGVzJYQ5wwdHpfam3rs83fJCOvpz3tuQ/W33Nnsy+p8Fg39WJwwLfYxdn49GorC+Hb
OniQpmAzXVMYfoyyQFk8j8ggoyExsF/lVsvtkOyBO3GF1GpBwAiH+0w1lRvnmdxGYXUdq1Z9WGk8
SyEDsbXVsQ8q00FyahYNoUoXFBAmxgiY48C0eN0UuLZ81Vo1LNt//33KdlKJlp5gxj3hAIqTzRG+
WPWRipxTAqaYvByXbw1CDnKPc4JVogL4oOByIhLX02rgOLiOTlMKs6P8Kr1+CB7GM90yXR80V6jD
VIkA4WEu70q0mDKsvE00OjaAfL3GRBtmMUjXUFXeHNIUcGSrkkPf0PyLHtAG/afk73AzE5UqRKXK
AwOref29ovHupTjKjKaek6vzhZeX7vUX1OljAJlYw+AoT4ndEscw6xMszG7vW9Ig7eT8mLBa9gbL
c5NyR3DqM5bztiYr8kLjY0tRyFdLG+wt6h1u1q7LQ8ANH4QKJjZM9e0vbwaT6Pw4sZ/djGsOiEAw
jh4jCS70gIAWd3NQhy+wQtR0iTcACrzIAWj+8ipLvDW0bv9LVzts21wSE7vzLwbKOaj852Id1OF0
yvO8ZBm69sX0iK2UqPHMI3q51J3Ju2TrTZMx/EPso82sarzVvbkQjLY+7P0JxiCwaPSXQbINj0lr
iPuywnhc0w0pNxWsTjZuUiNVbNVpPAl9+rUJA3yGxlePaAsaI3mcAGC77lD89m1EbOkp0C1QoXcC
vN53GtxEjHiYW/1tlKKW3XQs5SjiNux/+C8oGvEloWJv9jVK/R85HS9dMUz8SBhS5rMS1VY3k4T4
E+VBVq4zxeEXPbo/s3nBKraz6yN+XQAQ3qzDfAdH0mv2roqtqIA1Vb3DtsGBd77GVMAZaXfbBEyo
0L49J4/9rD3ytaLBEzbhG9Im4FR8ws5mLXsb3nxrEyTXNb6C1rTcpWVCNCHPIhffoT1Mjj2lXtEz
hHb3CEzwrywuOd1ZP4AtKhQNB7pxKv6uNgO2cJbpyrTDXY1wn20ba9M/4BAOheEgAPoqG2b/Do5X
VE8KgoxmWy4CZ/I6VdgnezmD6SNz5PFUzqlM6UqjJqIJOEn8BV1gDkLOSy1w2ZKwqu+HD1VxBrcJ
YoUV9d+w2MBIj5hN7HmsWN7Wf7UfdMQc0MUZrcABN5JqU/uBY3M3mxYRBY94uTUNFBqWbSp1rH4N
3HjQ+zpLtORm9IJJyQws9vF3sNVkRuYaUee5u/GgWfo4k9pdijkBHdIJ/dRLOAfwU4dzQBkrn06M
0zJGTNX0oZQTQriVeXM4OMHwX7aj/OnsXwYYdIYbaNgtCdJbI9FWklOzKtFYvrhirpMlZ08FVuzx
FVe6teiSrvGl7pWSf6YtHZq5vvJsMX6Z8BO/uPcxCF8Hon7elgIDD7MtBWVh28n/L9ugw7TZjtE4
729n8COBzMv2C54yrTniIHaOxCL+mOnac+G+Wc/nq0IdbWdw5kh5bpwIncLltAmUDx9ER5yauDvc
8+/Iwlh/RGr/kqAiL1KdXCwGCAD1eaIcmaBqZCYqxxyLOzOSQTvUFlx8oKRSGr/T908JOu06feBp
xSTUt7sksilTW9Wrk+sqyMrxAb3CLjQOIvd0bcgFfHGH2zIhOebGSTA3sd6SQvhnyZd3K1Jicin2
bmwHUxJL/WOgGhovweEcvnhPRCBa4gT0i3KKShwKHEYLhr2aLEBta4R0iRD6Wv/ZDAGwla3agpVq
OfvBFqdbiwAmKSO31D1otx36Gx4kCpxOB3eeMEfV7yN5+AqQQKzev8noF2PJhF4KLe/JwFzHI8O4
khCFUS9FMSWDfl+Zsm6/sMxkU/s9+p8l/92JfIStcP1W09iFLwByj3wf5IaYhGH8ropUdJ8+4iB+
0aZf+I9CInp6KY+onFxia1BVABLWXNi/N9PqD4lbVqsosdGhssiVHOJxvnC5jESJ36F//IqeV224
LXvZbphl3JVP7GlhJk+wTWmBFS6HAVHM3G5wlp8BwEfdW05hS4WkAguoAwjPGlK4Gfgufj/F3ZBj
/FmzKu5kcJM4VmJZsKcMXOEqtSJcQgIWroc9qqtoVQF9jSx5U6dNFL4mqEU0cJrXX1AuaBk0xlxS
sAWjfYCgOe5Q7WtDj6Sd/Wqjt//M3CJp3pI5DYu2YDvJUWOgRcQ5fV8WYauLufuJWSgZYXdju70P
prVvG3FSc0EsdDlt2lrwJ5DPsvWjRRUoEaRz7H+keDrCmcOrdu9MKKysnUHvBagl7WQaxC7CvBUl
sRF3RBi5bk6FY/LroDBV7iExTNjj0iRGHVd6wWhvvVrdBB0FioQhusNbU7aoXMVqseyntjpV/1yl
jgJJByf8E8tqVDvGqRSlBgabcyQFblagdSJlNKbDWv3lDyTmmnYs+Q3J/LBJPsAc3Rl+D6PVFlyF
lilFcCc59LH+sI7PyhL8SzIB+ihHle0I2PDilZiHa93QHIGBjlYke1EwMMliVw1bBUjRZQX71PBL
qMmf/OXUVxC/NAoB48BEvcBeDZSshOeFTxK6kcedu7EaFZnuLDAH2CkrTdKtEm5EXF6YowZassdY
jd8Ksd6yCQCdpEx2zIssw7UqGZAADYAayBuGqI1dyJiSTkgkZpjG0/BOD0LBXpo09sAB7jIgCFll
b1rE4zZrPnGiMZGhQGdm+3WN0x1cd5Jj3sZ1heXb9b50rY+1OKE07dOjzSxNCXvytu+JlCIDNLMU
WuE/XK/T367U8agylKvLmb1qoFdLIyvkTvvClZeaxKkA24RwlNHSqoejAOCd6XAvsDYE0gO8p3GF
kGij0PPHl27KAVFjYRgP9z2igj/93iDBG+P5fk40vptIyL+5j1rrK9rej0YUbLbQJBrxp/Q/Qebo
DQSKuT78fRgctpA1J2oztzb1ZiSAIReTi17ZefDkzQROFwnB1J7T+SDEf/c8Xk8KbiKdX0qR/e5E
qlxq6dK+m8NjneMKakXB56plAp2feFbMCA+gCdRL8MSvXtxePM6zH85BQjtTBJpr6/AYSWRI0hxC
NgW1jDd98FSF4koSzj8fMPbRmSFXRba9fUijNQm64yeP4L8Y/4gE1KIwviXBAVToJAIZCnrFwawk
uarS7PEmbH8WNEL2POZrskKeMyzzAnA9uU92riMC4Sd93wD8S90G0woHfcerWlhaBfgSJ60oImTr
9SA+sSJXdNBl50OFhmOmMlJWNxjSVVA160stvUzkRKoWyOvykuTOVo/T27sgHn8a2Ff4x5gmbKoz
qJTOgrAoNLxN8pmcBZT4G37pMz86f+n9bvUqqnyeoyEaRM/FxAWAUEkA7ZtS/XRBIvDYhg5EPBUj
vdhiJOD4enl08CTKtxsV59TZl0EhA/iS/rm+GfVRFk28O70sas4gVGPEw2027mchhyL3dggYIEJQ
xA2LV6tq4ZJ3Btlhmk5L7DOshYCUwjVYI+kvkrXsEW7023id5x3l/LRkUSWBrKbfdy7dyrzTpY3l
VTQGCRSJ+Yo5drfKNeZBbnfs1ssVcpUSDF6l2AxEDzfJCsHpO+/t4maTWnXOUl5VKtKk7CYuOjxe
o2qEIBiy6u8AjIHG/A6GRg8WhDwVtCWsuj7QQMmMQ486B8Of0iIfCb8RE6p2IW2wY+mb1bRQBG98
oZ9bg+bW4TR1enIhxwmURtLIWOefZfTWtAnt7PR9QDgmx4ywPA+J0CIpGoRJTNWV9KpEdGNqK7nx
8+07U9S/mUtgX1jvN6EVb4R/dXAQD1Yzt4xv1mSBioC+Tr67/TBS1ktljR0WvHBhXF2pkeY9UYxe
QPtZQwTz6FI6BP7x0V1ky9rA1NX2aUTMhaisF5hu6UoU2SPE7kbi65IWVFCwposX175Evk6tewSz
ZdIF/rYHSqkXN3jZjFUxLR/44caqoFeBZaF9Hj3eDr1SZYbNmu9k6jCwFmSEhzu4g1A/3LUXocJh
uWye0hfBV14OI1b4W2iVlvvi9MV+5oT+1oOGvlGVwgQo21AmhwYyD7HXS7oW4ih/yVRxH3fcjz4d
AqR9ZHgpptsrblraCPV4/q2ClSm7l7kDOvjhGod1/SYhsrD19xktDS66TGr7MzQHVcK1EujQhUC6
CT/ivTB/1QLJlLcd4GIClWBap9MMAhzuP9LkLkMLmhN08h00NOJW7xXQgNSaanqCETcKCT1HVIPi
ETpn9yMhS6CPhJxmDeDG14PNpjJD9jIZIgdbj3Zr49q0XcBNMmliLVjR5P5xG365SlplqEtKS4yv
U06/7Jqd+Pnnt3wcOizN9x1XFuiWZjqRhJi4dM4YGCCkfNjOHNjcD1oq9/AgtsGKZzi+ndj+KNZR
tfFU3U1ZIJzlg0Jno6WHSS0GL8VAaxRzfP2/UjOnq/ZMGfILXLZhL/XETBX4iUXQEVWSe//G9++c
MPMm8VEChEdwKJ1RbZ2hrYJ/urRTnbnzG35owXUC1fhNtFwr2aUBUj/aq9ixjiq2srzlOCwPFzZv
GyZApjWceVBUwG7BxK9wj/YhbIFKFcCOXAHjiJxjsQkWB9ihfUYdiKWV1KZBog+pzqcucDTeQPOb
NhZh6GfjQhcFTObqLzzJkn0uBDe7SJ/2S7NJX1Eb+bDG5y8xutd4RIEcNzvh9EFz5GYgyXtcWFic
puXIhKDsJyWXt0pfYu6rRQn95Tms3oOg7Ned1AnsAUm0t1wc2acIJzxVpBDFT1qtEtmsqXOYrVhA
/CxTNwy2MyDC4MgXpywQa+bDD1imzBRI2gPnwtafQsccG4RMQ09WKM3J9zs5PAFF8keG7X8FhktL
Ax2NyDybVAZ0nn7IJIqGbQ1w4zQG9em4iaj4F/1RrFCbhlEz3bWNLKcYg3Wg4tMAEX+uTR+B+BgT
OTiXu99QMYQymY5LAtr5VI+c3/ECvKwc8G6Vn9tBlRS7D9Qfp4Tziv6RqoevNU01XXnFMVaSYEh7
VL4L23yRgZAtHzqvoJ6Q2GzoQsk0Dd+nZO2u871edUxDLvN7Jq5FpEbV8a+LKcTf4oV0Uu9OHk7U
Kk+HcPjJA7bYpbloCNFemj+4AMziuzXlCTPTUktyqCHqkOZh8W/Uyq244B6LwN4k3tzEOWN8wHQS
ewdRP+UGzkvZmnLc9cmNY4VvOL6rRWaggK0gls4FURSEep9V5MGmXcdyqX9vEKDXTlOiOMQka0Vy
TO4UHkFkTEvRkHDmsA3FFQgYhYc5UA6vk2XIVXQK/thZg/qttDBMFSfh0ubr4Fo0IwxGvaTPdd6x
0CJXhG6AAGX9TlWo1+Oqk/6BVkXXICdMEkZfYfLlNqcIaxdCe42xp6u2xpBG1rEdNDaUi33F/qrb
zLWvCeuauz+257kf1KOc6jPj/iLHjVpdZ3lhU2lA2HKQWpCBkOXv1mhGl2YmsDiixoxJM/hZ5SRH
V8fxYHmAkW+oR9ebLfYeWv9JYaj8r6EIsUQ01ZLmiFRRZJ4IELssKkYT5bnFCecOQyHSrS7mtYd9
0FhbGM0CQN0M6gPrWC3uIF+efpeNLMosyJ+HruX0zQ78HTdTtmej1yN1rUAjv7+XHo3uf/aloDrl
hx0t8nxU1O73EgFtune3P7qk8MKnFUQxg5ZtlIN7FeQhSRNBPzGMLPsXf/Jz9nnBOsaL6fU8hV1v
LUycGWVoxZklWKmHLpaDEzoqi2+jRV7A1MJwK6b6vr95OEgBPVpwdmMT1yeBh3MHTku7TEkcBz/c
Ybm1Tt7tmOQ/ch9rEq8DrH2gPXTJhWBow9Vnmb7JpawXSz80f9O075m4XUikX0u698DfCC02NYeP
wpRIxVJ6S0HOhZ79Ihli/jvEVwaxM15/K4jtsQ9n+R0ehMm0JI7c90g/R74igPoUSgAYl+mElIJU
Y0aj/g/QVFZEm6ESRvRGixtzwZfnkTxcy6nJkwBC5FiZ/yCBKDBv43mE5rM+/6n6jQltzz0g2Cr9
RtHQoDNiuqdPtGj2LB82D9Ts3VtuYG0qrdxZGOBpu/IMjagBsITcs9+DsbFYqb2OCpR9ILCKPGgM
enotnqeYQ6QDd+RboRJ6YKVtYlMiUEZnI4CPgggforzXU1I/Wr8NenM7e3Ya64aGeQOm0TMgEZdW
kIC/yUKwxEBIqkF5lmNmb6DlPBqJv5GWKjsBLFBttmTOF944WKefWN2fUKUtHqwar7oeU8d/jhZh
+CN3OJNLWsLtRHcQYNfHrUgeVs4CGw8+k2c++Gq8UD0DONTSJMYgz+1qcKuLOQmZc9my/EwyZSVR
dINpeBs+3aNJZkTrgBVrWwRROaQB+EiaHqi6aI0onGCDVi/bimySWDiL0NY4Vf22hDXW4S8SxRMW
JRI0hNaOMUas5lrhgUXoyHuaN7aFY6gw7ZmIIrHDDoojRme/E1WQI7oPXLqUvZhGtQaf6siPP6BV
MU+2YZ10ROFURP7DqHO935qLXh/v4RlwmKCouvjKlC+sawRiJ/RMFLk7x6hqzPZnQsyMge/ShBmo
NX+IlETkN9SQpg9UK/yR/nQV3mUUx+I8zuCpGt9hd2HqUtboKrkuHWbJcXKrgWCT3YwguITY9Msy
g4lMpDKTA4jCKHIloa5R61r3wZkRJf4MC3Zs/NQKu+WXefpPsua9ew4VoZa+ts54qgSmMNRqszLj
oLdzFzqM4ceT7ADvxuKdsyCjfBWtnqeXdqrw39u4AisOPRX8EagpYzgv4S7mfDzxtTUnOTFS1bSY
AD23qnQo86dwnVpFJxeqFl778nJfxsUP2aefTh/b8afHcMr243LBiLxTSfaHeT49vtOgyFNwE/Vs
a3jlijPTYk1E6IkD1eG52+KHwW+KvuOAEVu+bpuRpx/VE1PpZYdeDOjQmmaLEJ0qtzLHcs8173w0
cQStUNqbD8LGrVQ79B2E5EHxdG+cmPaelTL+5vuFw97t6Iw8vegqAgGus3wP/IJIB8im1D6V5wil
QcFFM3kwQ56vxEGr5zdTLiVoWT5e5SkmPGlnIO4FHGat971qExtrbrkjZQ2GMNxhu5vr8KgWnXDJ
hoU+csbS2UOmcfaho0Zq7WKuKjCrhfsuFNxvLu13iJnLXtjsZrG4yXNxVqESsn2c0Fude947S/bp
+khxkathq5MMnLb+ij3Nnp+yAy/W3p0pmUG/1r4bPbI3bPEKZLWEy4Xg1NlFv8f3g9HiDSaWpj4z
xwUjYi6fbdkFBih/h2D2kVh5l5RNCFszmZURTJbDhWKI1KJkXZ48C5W2oJW+3aRqyLcaYolevVdB
0rFoZVkqvd9a11jLE36hlij/BtjARWl+HMQheebdbSnC1S8X524r9uypuW1OsaH0O4U6uWozyh2f
QX6G7kEnWaAPxWZeH0z1IVOA44s82ecEuUACEW+0nVpn0pnQQO1sAfWEdmFfPJnqMQzqEvyqQEnR
FVYUIZRzkUZqQrhtm1g2Y+ltDzys2cyoNzXquWYU3CoV03O/KbEa+Vcj1+A+NZ71VItZ0D+sf5eA
0Nv44jXKFSv7b1McjeRfC2yIu/mfkE8f19ltt7Eb9fcy4ENDqUmnvvrD6OgLUACL5ucyfckER5gw
1SuB9zRFznO9SkTX/sIo3zSVFPyFkfatBciG6avHHYZiwrznoXjbCMXZ0Dq8DkNNpMkSZE4Us7I+
XD5IOB5+mej3wBB0OQBn7IT1TMLaEgxv1j/KWEXdo8smAsX0kxrXn8FhtxrIQhGvpZWqW+lBI2Gs
OYIb94Xy/vr4+jByJY2BdbB0X/4IiyuZ7Rby5ETzyyLJWDPZHPYY1f7csivevVtxnPuTixyFbjvQ
UTFq+Q5gAMQryFyrV5/A2msZQtTkTjR3QU8TNpk4VB7yfCbZQlnAcKJJkjAUmTT6V0JFQfk6DuYz
AuzL3KjApQiNUlmiZ+y9NZ2OhAoaFn1O3FGZsKOM1fgc/3DipdMyyc8fZbVvIZmAETvatJnKqCFP
xCOu+PV6UHsmjTWzjYPyeg4Bgt78+/5z/Du/32yBDu0aQvQLinhV13PzLDz1zjC68cFHsArFGbXH
bANao2+EFRsHPhGv4PvMWUh/jXcVLMW6IB6a4Wtm4W/LUAur1I78dq9+gwV41po2b4ryqMcn1uTZ
WEHYXbAi0ZoeLcPAnx0Z9WBHSPQ6PWtpVP2apnrnAPkWl5Se7jq0W0FszgpT3r7HgFeHHckA+KXM
5EbYvzfrGRCd7M4nPFMaAHWpGxNOVWYRw4/or88v3cHDI8xLIeISR0Q70AVQ9cXrymB/m3pzu86k
9KRiu5R6e43KsfL6BZKfvAO4VFpRERiKlnQayCwnTnQx46PeiPRe5GENlL5499PoYuQ+APSAl5zh
fJ1K85Ch4eIiSIDds6jYv+sVjSl2FlucB+CkyT2F4wYXl87zSPr1mJYB1Qq7MJ5fBvBXjA/03BK5
go816Ih2bX8nS8iX2vq1LBs93ZWCc5E24hoeuQEEMsLCEfmghCcmGhDJZWpvzR+y04BptfT9oNMS
hjsOHJOhrLj+v9Qy/ylZIKf4pDT8CUDfuhe547um23GhNDjMqSY6oKOcPn21MaZbVNmAUS86DfCt
K0a/ARNf3dTYqNZOQU/dSaopIVwDrf8GlbeOkuVeekh3uQuwv1xKA3X2i7Zn0JscjkBS0wrOJAG6
mQwxibk3/VhSlyPPLFafmGGC3hMRJdzhzCaBVJ/1tAre+hzcTj4oco9DghP+9iK1aN1IoibVC/o9
kvZO1I+2Hsvm7kvGoGAZLsC/ENlOE6A67pv/mx0Y+paSIud9m/ynQA+qw4ax/DyMqDj1ey9Po6/k
zNgDOGae/5HLq8Yxw6TyBO3ZLhgi3om6tRUQLSPgWH219V51DnhD52XAC0obnfrOIHgHy0SlnGoA
WDuU/v/8EFd7HxKuQsqqDw01UypYhg3hsN+QKee+wnaDjvpA/u/6kQoPq5Rk7oKPZ4OOFvONYT0J
r+PZeV4TPGZv7MQbxQINIXfMuq/vV7vDo2e78ds6TrOajLhMQOrtTT+DMotk+ksFF7wTqNpLWAj3
fjc5Ywjbosu/9+it5cVo59btJRFDbuAH8Kf4134ZRVUxmThkiK7Q+MPXI26CCU/VQb3DUozPccnk
N12iYCqDEoUUvg+3mAZBFDX0aezK4RpfriQx+JFqiaI0QTPr6Wvxqcg1uH1p+HaNnDA34etoIpG9
qhdnSGc3XS3WgD+7kESUKLgHu75Adkv7HGhlXhOXvMcvMJepbwHQ+IuM+8YmzldBC0wN7bf6MLT2
g8KXcI/hItEqmFW23LXwvUyV16dDQhIOD/Zz9+tN+DB4niqqnfQIlPDTrC0mkL4SDQ4X365UqndD
G6bU/YPMm6NjbY0xLR3brMzP5ETO6NSJEGmR7WBn31lPNwUqEMSCb30VLnu0h5zk5MUZI0f+S/vQ
z24D+nkYPUPvuSiXWSKsta3Wj0SHDknqRE7pMVfvSfAvfnihTdlS9687HFeIeaGAv6R+6SwsexMq
s9FBumkKJ4vqyDHvitQOD/70hnJJKzuxbLy5ibVGd8i8bnHXeF/Y+QhJAuttRXZ0KYzFY0yMzW6l
/XcUq1ux+G31fV4POQWCIRpB1VvL4g8bd5/HCOuOYJDLEkfcVp8xRMofYTgtvSJ4lL+O8bLbDH0m
B+6lyk2Q4FkktnGwWzbtuq4akbNWwHveotGv/91kPBqdAFHjbzk2Z4han2d7COtW+dmGOzPTR00E
O8UQFaDz8Lk7dEvizeuzYqiN4CNBwNuqCBquIq1uM4JRGLF2w1XJiMFKl4LsPpkG6reTX4NYg/Nr
p8f3QzA/oK9j68LG3fM44dk1tGP64uMEY0L9GLLU3ZV7a6Sof5a/7gh7d34Mx9XwHkJcRIxz0U26
7ou84BnSOZapCMYd6vHXz1WCS0/pvLm5ZqQyFQSLwfdL9tR8CrOMfRF+QIZM7t7gTBeFoqcZXOWh
5E3sGrDlxoFb7sHySglru+Z4H6bbBxlTjt4KIc147PJsVNqiJn3Kmw6RUs2wcPENdnG4r3cDrjvA
O3h+VyjD0mXgQ1pFFhcuLx+6GZRoGKr5HlyAQtKzEuIzS9578BhnNuzX8ng55Hob7Ja1tCsOqIKO
WOP6a97eBGKyWNF+gYoEXtUkGO9Nk9ZjgeQq5murniJHVRgbnTdsjtN7HPG9OPndlIkIEWHxBOLf
WL47jFb2J+lP/JTFzTmy7sMHQ/fjvVkaG+Lmg8MZnzCkMs6fqif0QCt8QDB+JRc0EYzvf2sxD+xv
3XO5Cu7j8NgWU9isxEwtpkmeNL0XPYsD3pV6WqCgsWH+YqzskyLIzGzbIj7AvYBuM3K148II2HDW
6M9EmVWob8HidKNRvFDi3akmsE8DvEOQnaaEEqk7SKJTczrAEmNIktbLl2l3EaiWLWSJsZDASevX
vg5J6sJfqQMe/mqPxwi3Yipm6NBhTO5X5fwh29uF6VOCl7L8JXzTnkBztTdObYwKqk5heDB1w9fe
LzZEBGVvnhl3JF7TEA1uoXzNNmdlElxcvFj/Sn/3cAczDrBvaL5G6fn5TCsNaUa5LkiqR0Vl+mHU
NNHATxLtGKWVUMk2C1hV74whsxos0ArJE7FHToj8N41HB0NyyEn6EIVx4nz6n3y/8SvIxzqWtnr6
+EhPBNqtO4Z15zx1+mtNSUOedwW2gPGusmBbPqVLgHVb42x7SoCkqNbvcaeF+pr3hb+wH9sxVs6t
PFjGP7JkIiOpWAS1Ks9GDCUHNKwVtOv20x1+V/9giAiJ7zr1z4N6bC42fgObEu48O8JFjlWfyjqh
bT9mYNvP+Klg3wJyVshCZqnVk+BJv2SNPgW2+q7T/tJizUdSL4VqAUdi1ERdg3R0qj0GAjXXLNpI
vKftH/caJJhX04D7dkFv8Epahg/Ple62adIOcqj68UkWIvNAjLFNgIrxrV4/59qH/GDUcoR/Mg2w
0KzaoAm3uj0GbXYf9/lZ4vr7x7+TwF5ZLvJXRYEiAgimTB5roYnCqI3v0v5A85LknXzx4S3r5cCR
px4mPh0Xr3BCXRbIyI5dp6XL2ZXskfIzZagkTeKOIMMno2NMOwIWFSA68wVcrgFFTuR/D9ci0+OA
V4Wev6C7PzbQ6nkWUiib7A+ZaOxmZSteg2BA7CA/s4GrqKuTaoKfKIKUt0Oubzs6Y2kfMBNmtIfL
NgM+G3WncxlJGzxrDP1qd8CzCW+OAj04wh4ANdQmrFcl7qJSMB9OvtdRnLeUT1W6g8YCTfUHfRYf
B3h1OME2QEErVnnTRig/OVwIQy71+Yoc/lp81iQymGo5eVmfGxXCGbocT1TMbnEiD9BUOWtUUpaX
86FeKaq4NQyYwRFeFCFWUx6oflOIRNx/EC4Y2Uf7qGHQdKJlXOwbd2RiraUp4PxSQO4Z7OXMTtZR
JiO3MUtxQd4jgWLCjId6sfwllqVCOlnAL89GWmPp4A4UEx1JGS51XLHRf8THkhWUH+tNUVZO3ep6
R5ZXM1dld42PL4jhgsOtQLfbmmBsE0PHXZeXZ2/PGBvC7oK5P+dubf+78zr9VxOJRvUCpZFmqxGc
6rfKII0Aw0Lx0STNoJojXf/IkomUkP05/KbMciktYFC4iFcznWHsBu2iu0p4GVYbnuRBYDcQhbn9
644H08n3E6US7+PF2+ZGC7XVD8hzN3TEFDEU8385DsCzP3G0P8TLJ/ey5Glc/y+7uP8ZAAr0s/4a
ePyGTQOh54kohoTvk9FM2gDFDP+eq+f2lohKb1UHz0mK5wf/lsyEToEiuw3MFfp5nYkEnm02+xn8
SUFetcSpOGxYXOskF9R0HsE2G1g6fCQZDY+26kd/XBvsYcLxXxShUWWLoDNiDlfyKuZD1qAlzCX2
ziSp4xy5dEgGZTdEQflwtlNuJJHasCs5ykXQlLt4HVV5NFZDjh32UI+bco1thq6wJRf5t0jXI4KQ
HVNoddUIKnn+gyr0sd1rrvY1+4vrpXbkUo1RT/g2vKbIa+xp6Ky087zWi4R7PB85TfMZUd36n2nv
yF6Jf38O74xNHHCHt2Hnp5vKM8qOhHh9iyA/rt7vvDJC+SmCaJQuGClFVe0QuM+OwBMEwQZBEnxV
mrqiuYSVsHKocahLF6rXQD/zC+1ezETPvOMwbCbjV5Kte7LI8GdwPNEf+sO4svc7muvE9pJ58KWS
LcTkYQEj5/ysoh6VJLsBtmsUBqzjaHU1+ifHiQiy0KlLOlfwXNXqEpVfsdtCmNxg8Olch/vP2t7Z
rTNfncbMk8AUeLz7Y4EbX3PGR5BC3vP2Kzck/s0DXkDkaBY4DV7u/Uz2kmpl0Ps89fS3/xDiloDA
M8IPvV9VOQrkxc4H0RKbpwZ/oeaKIax1yHkVJ+83i5UhBZKRdfTk55/L1wKOHXoYER8I8cde6W6F
sylY5ZlYi+Pyo/ctiXK0e//v+X0vSU6TRlNdSR5xx3tP2toh/XDrZBKHTtAJvHghWySLW7D75tx8
DHdeVCnuzDcZHNUyvmjUcDV2VA1AJN57xmM56h1rFfxrztfN+BBL2Ww8yQTw+iATKLrcuGZWqgpr
xunjB+Ui/oPZ3FN5dM3BXElTKrhzjYCbJgHo1FNwaldhcIfAaNinHx20gymEx8ktqrMNukypsUVN
rlRqhfwW8mHPqumnOj4lNddnrzQcRquxMPRr8uWeNkWvf1YKisoPU9aGXFbifeTUQZQ4wP7o/5AG
6SrwmhRCTt0sVSV7BPBblY8uvF0ySBWUSvC3bR/xrcIPf2amUn8lJNZ60NCjNi/+MYhr1azBVbM/
hBHzu2ghMdTl+EbsTwdeHDkHDMiUSal99HC9py2Xln5DJpSTxcIxhvfgNES39Kxl7w1aqYEAayWD
JUePTq1pYlk66zSa0kSzZ6bY3n9933gMAY3w5CHprzJJsuo50E5QHIarh/3n4zws6N7BUvepQDiz
4wzzgOdIzFG06u639inlLf9w1MwyMDwt6YIkVA0jUVEMeVxDoPhbS/mjWQrHNczxxDP3AjWr7SAV
4Q3SH8U9f1aleeAm3+55Gd3UfokouVNrk8vLvQQJJJ6Wsx7sNiY11PMR8Ixh4TjRf10W7Y7mE5ee
Sg/TJzhn9Km41M42FBmSEZjR6D2OBoW2tzpx4SFgQHcLljR0qXAEt2vySnRn5F7KYuhCCr5TPzL2
rGJGGsFQl031mzcN118k8ntw3hVPNgebsI/OyC5jouSQr7Q12OfzMA5MarSpMd6S0cB56NcZ1/w/
UYwVxCu70jVtkp5ezNkU9xTigbChYrIw1/gaGJIpGpTe5y+ePYN1ND0KclbMQ83NqOgGY7R2HZGs
BCOrmmu8QprF4/FU9+7lPokDwVjzF8z1qUDkKo7bCpsFs/Ky8Cfrb054i2E5PB83VSjmFkYGjub9
RKmcBWPi3+2G6HFMCxQjCyAPWNNDFmPkSwMyrpwMM1dXgY6yxT829QrvlSTSZBH6JbbOwuh9JhSz
bBaUSjObnoIpkIsqTRew9JoggypHS/5PQpHYHh+FEfwhJiy0TdWnnE4sfIrMFNSz5JRrs3chEuDT
4+/8wWlTRpWE0Wwz2VDc96B1AeVKN0qCZyFoslECsjMYu8Qnao79H/Sm9AYF2WDav2w6hgmn23kL
C4nYqtxcPBixAdgrJX46nxkMpH8lRyGRx0E9WBh+pMQYtyFqEr0V3m3lSvK76VQ6KeFUak62uGCy
s+zCiFXhsUlFMF2RtNFDPRZFKLAd30rhMkeyT4+gZ+CkmEepr8gUlWR4KDLuen9gI/dsrfR/h8Gj
Vdl3eQZRtTi7he6WXxF/rtQCq+XQr23ejfDVN2oPKORhq1dKkmTKCkhUgaQRB6ETCq4UyYF86+HB
+l0BKWs0dhkuW+GjsPl38Jv3blqT/Rtnjp/OzBZ3CBnQ8BI+ndAsF3bYcrqy3Qf3XHPhV98ds4C6
Q49VlOCy6KGQbqUpCQRZmy2f/0yCbYq3Hrhw3ANok8siEhe8v3P91CAEMuswkBPj6jjXM+7mcE4X
vBoVWe11UWTfEP+tzcH+qpPyNLzIGK9If5HysnEmOJDWqxl9rUBj49wGGlL+nE+08W1HuyLoHU4W
FukWJU+47ltbjDcWVOLnYNk6FL2Ky4NIGlrafNuIZEshh9ts+uKAE6zHDK5aYQtFnFhxX7YGmhjF
Dk68AVKF8RUaLjVIQ9gGOT3cg07GNhyfUndzkvihN/qOUncsA1FyGlIZfLGGVYV3sqF6wEswfi7m
xNtfUkFn9p/sTD+IVbkJbmi7+jnnKxx6FiVnd5g+IkcsLy+HxfJKkeko4JWa0ttxqfotTJMGAO+C
ftqxDOqy4arl6jl3Cwwq5neuPZ+I8ll1jHR24EtioFx4yxUKfSo4qi4cCJe43rZKUP6B15d3VcIO
2lN0q8h9XfMKyjtP+fri45vIaDTar8MpN6lYkW3OK43GZ+ASg5/05X19OXf1YqfJNu78o6gX/lsb
yAO3UMEg/jqfDGXeCawhoXUa/qStHi1Asmf8cjndKRAyV/PLsYESOlrQWv9H9vqgObVutZv1sFs7
fh/iW/w7fHyDXJuPeDwR1dSSVQiV66zKmeE2Gya8MhT8X6dhvgZHNOoaLXY8NACgNMz40m/J7ey5
lX/J8r5ngAlXonZxY+q1RUQx5oWWmQhgU8xdsaOm0RYLDpp73VW6vqivNRKnRy2DlCW7+KfPdTds
oAPJ81Zyq+yVcpVQqqVprUohaj0AXkzSbDxhzTWE9evd1IREVFzuWlyjL/w2g/JZrqM1cR/Aswio
Yv03jl76v4GObNWGIYjla4unCL7k42Qms7eEw6B+QgsoYVZBFSRnq8QwXLs6TVcez2JuxG1jMhKD
Hgm5T0SPYegUXbzd8u0bk4TleRrE5yAJTMw8kRnlYo58oNzF2GGVtIjbff2fNqOaz1kxHYmYWQen
+rGd8dJ55q6IuINNXW7KQnWzrQ1BjLiLh1JgxuYQEYgL6PX9vUIxBGevWQQ8aDZ2ivfkqGfOGeni
gaqTb/5LnvqYYh8+WpK4u5HHzpwWEl1KCqd2y4Rf4fCUPH5T7c5gbIqbq0mQ8aJ4qs4aMlm1m9Fb
EzFQLHHrQDj0k7hWZMF3VXb44CS16io/UHn/cf9sp/9m75aRQ9Yk5xa8IB2qw65lP/pN+uHF7NCz
anSZ0ufRQgeA7ZIVMcLZXreOLyHigRjL0PXaDbOmwPwKqDcFr8wR5i4bcttLMy646eO6a2FWtEww
YbCMe6eDPwfMEzm2OkCHLbyTnxVMfWTCD3ndDGLBko/uQzBjMYtMpl4jD8IreLum1yfEBjHun1R3
pKs25JnSW4Z5ffU6Ax5Zz133DTzXz7exGgc90JAucKcYgRU4U3ZjIxYmAGiYazgvzt9GqRc0VU2p
G5v9ErbkyBcnHCtIsQVBN3b6zS3N6DJsvB+QTMu5ifuFS9fCCuV1F12XqIBBnbUYiWGb+kxru1HX
cGjJCc5BA9tVY9G3fal9aTHikJZGgSN0clL0e3T0HoNEOeZv1wwMFmk88rYw4AtE5ZGgUDEZtjGL
NSeVV4zMMnYZDFIETVlQnu/unmrZBxNROiWfD0c/oGu1RNfIZ1Cerz3iPcdOVbX7IhjZxuzoRMCj
1wzrQs5c1tg4ltiB3FeEBt/49iLAtMn0aOI+/cH7o8qFo+BUFcKXdfFiKUZDuhMlSWEJg+P8Wbfy
NZl8fDkiHRH/f0RmgjNLu4PMQdqLdc+3Qtt431P52u3IGwxlMIw52WMq518gAVHpC1e/6RFMDGMS
o72Yg9P4a48AjYbv2VWXhVgepPiMdw3XetvbLYZmikkAtpLUCOEosqTvs+g9qpMjscUH/VZpEw5W
qPp0Dggeluo9fELgatc8ke4vIhnFQTj8vcMtYipX+O+Cr1eZlDcp9AV+eO3Ssl4qHjQciFM3Zf2+
amke7rj6gC1lG7apHjw64ciiO48A6E1/x55Mg/qtHETZ0xGo759m6oLP4ClQgEi18w+KBXieiJMi
FxZt859f6HctRjwXB1OpZxRzAXdpICXkKq0H+LAZnuaKGUxdF0vfZKxu0WeD9zCoWC8teXXocI78
CUQBeliFEHA6/ntmJFAbVOCEz+FxkrZy+VmM6ZIGJtGhdf9eU8w285pRzEq0ATjEV58F+BU++Czg
0lJiXhbGnLSYWb2Y5w3fMFhQh2nyA3afs6AaF8m5So6BjGNvB0UgF09I5Sl/gutillBU0yhjPY2Z
SHp5fHdFLZOgAHYqH2wDJykSEwPxZAne86do5mNxaJXoiPvNRJTDEg+wN7KgmztsRxdT6Duy3izi
OA1yX7zIP2tSofhvJscm9+fDVrzoRQ6sm9u/aPz9DxEmxxXMLBDLn/jJtOxJKegVfhPG7BvV0way
rM2zhGCiFlbO+4LbQkSk5P3dcQ8ncaKIoGVyoRcduYr8R9dDHP24S0hpwAehmidpivulh9BthE+D
Pk1fE3AfcJ1+NEPgX27+EJ7SmLKXVekRo9IBqYA2GAR7V4ifmUQGdbVRh2fgY0HX/gO3IXMn9clj
hH7jYeMbWccQhwhH8vfKKy9cLcolZ1nK5GvREc2Wrq4tVoDGjUUeLJZqZsMrG7iDCab0OSEKbWq/
tdrIM8W5y6C7jEbVvD4YP5l4ZOCiVJOHK2rX34lzuOTIqNIWcWSigrXYVDHh3lAdj8DHU7338UL8
qUABpLRCuQUme8OBBjwSNvlkdl+W0mVmkX3NYxrMMCyYlSdDPEEwD2PXDsVQfPaquncXw1vUKdjE
THjkyBEi6QVRCHtv8Bur8tRaZ+RBsjc9DF73rVOg1YK3VNo9leqHQHryq18+uZgFRnM98c5ZmruP
ZAc55WsYeP0qm1mEUU3hLTRooj2Wmczk1V+8+TAFbzrDtW70JGFj+UXsUeAgg53X5IMMCePuDc8d
2XUBQpjkVF1ge1TY9hCywkxD1xuXt5033WzOAouWoQF2z/0STciYqNMtSwHLerS7Q0vNarb54/dT
vyuv/rxJysTo1KCqubKSeI53uteDyfGyIl5ITwwOx0VDjCQxBe8Va/U9zg3g+D3D1ru8mYGGoGPu
J00p52QjOlbIQD9ZuBjnJiZNQB62RqFWGLBXT8gyEXO7L0ghuuir2hbvnd5qcJ2f2N0lbhDPlB7S
OPJ79vcSJdshB9PgtuT7lr/zN+PKLkBcbPuPtGYVaklpCjJWOZtYOO3VsMe164RNj94XRdWc/EWU
vKqSyItbGCgkanjWrTEBm7TtvwBb/AVMm1OSsryCnHlIHA9jyt8fZX8p3/Qn3K9K+O9F8y+jvXpq
2BLu2aA8M4+/IL9lk9QQpwPSJBRvZUpaAjozlyyYbd7xiDkgE79y8rkBtEt/yzcs9Dx+1/NPN7jC
sYFkitw2ukWMcILr3sZJKqf3FXDDmvVof1djc3F0ZnWEkn/KDbFX9e64qIDMr5lRlq7kJ1eVb0rj
sfoNCpuqwpIkuufuIYOQXtrzt9aa8l9bLVbdfeis8gWW554yXz0qg0+orNY49elerNh9DDTheuQn
UPPQYTlwrOFiE6n0X57DQb4WQL6/anYvBWiixd9VX5i0/dP0M8KjMUWo+FVY+A0dowdv98i9EnFi
Yuy4BtewD0iWr47anV3kWUhGznYfabIco+1CavHmE1zeESvtDQWvsugV/x6i+538bFNU73hcQhvf
YDVj6WDkyT67KS0pECgN2CawKqiF3I1BWcpEf3uzpeEL7yRmUftAa9EsmXUynetQlDxvfZi/gcvs
W694fHx2VBiNOxNd5s5cD5Hi/AgFE2FgjDG4rNYr71k7e8fZj7Kp6ChSXIz2td0qjHLuqWWaX8Cl
YcKCkcIEC/1Kzz4+rNMr7M+LP2dd4uxybiQiinRgoVHbuYO+tQEA7rDbP31sHDB9nUktu2nd/M9n
exCVbYmExRfzyI1Z2hdmWwS4rcoIFRmW/7SMB/FQAkJSqsM6aad1zXJnKoyUXVVYq7fboG14wHaN
dgaComyLJXZhyOhxuXuhArhkwhO/SNYXvKFarFSpAeqP+BkSMX0X6Ck1Q6R5ZJr8WZzFfRid4T1k
/aumwt71yOacDOe0/BN9K6JrXuvU0KabS9DPj7d+zb9K44C6w3qkJJsRxqieulT2AuO7pIKnlJY1
/6cGdPC95f+M1fcCcJAqELTWDUcefFN8GxydmAGipF0QY8Tr1DIl+w8uzt7n5p+5qMeiBTqAFg1S
gN+z+cH19b78+0c8CHBlhGaxhMOpeHwWS4/sqtFwzlLRQ3CfuUawSeLs2NuSf8zuGJt/JoaMINb7
8r3ywahMO/kTzqWXLchfkMP/BXwvjnorR3QDE21qXnZN+KQFL8niBDU3tRa7Px1YzZOf9D2BXZXb
itfnu3fjUXvGfi5YjIriZopYeClz9K7YclkfGFasiWoGjklaet3VEYhfprdZOQi5FHYW/FDe0zqP
P2RrwfV4edbbsk7bjRAQPh/s27+gQ4CFOuaUHF9jNciHzv18jibAcYcOqIPrFUbd+RGM4aDWTG6R
2SLqCc0jEnZICwPVfslTCBMnJ9i+Rq29/eA3muCv4+K5BbvSzUI50SBnyZMNhQV01eFHzcsuTyQq
KF5q+WrNQn8IuP+IpP7q8bjkKaMn2+ZLb8Y4fIy/No2g25iKRFss/0ya7xd2B7kr1c85IDxbC2Pc
zBMUvS7rc7znMvt3bkIkctUlfshQTgrwpq5CqYHEiqxtAXtiVnp8E2TOSfpXEwVnu6PW5nuRd/qn
4ouFqGhQedqm//vtQ/iK8g5p273MhOfl9RAUJN4k0PBdiF2oQFB522IxNazsAsFLeHE5cJEFK1HI
+r+SWl0EmsKydyHbRcj/zeud6Mq7+qAKusnevFzP3w2l6JzSXy6vIOhNFNxKEDjGiPj9nmJKHQXg
njeMI4+x5QW+hJxrKxbwGTytCsREoy6JaRh16ASu6u59USkCmq8rQ21k40qVL3nWCL6GOl4QqYPf
cU9AWqkPyz0asDn0aPtaxtnNW5z8A8xUT4Swa7us0dOvE4WBDAtS6IjPKK0gBUVRBfSOtHwxkjA4
MUaB9N+3gIZGXDK8EEtPGPvdMlQ1ASHCZ3wLkjErKR2846ZSwqONW/aIfiLZdLAeqmjgAbcSFHs/
aFg6eoh5Rpoc18LizZ64kulMxMsTufvQlAfZOwpwPk/zIvhKRGHQhDQnQAUe0xVZPBvacptCq/VS
JfdXG8y+aIHXE7LOGDQBQL0fbABhyhdcD8GAjxepOWZ9aalcDkb3jm/+BxfWrIgt3jKkY0qUeIG0
zNFhY97FEv+N99JktYUo3Gi4+rzEQECgqpaYKOdqvkRl2yM9iFelzVNmsbxonqUMW3nfEJpJk60/
3V/Vz9sb5epznMrWRWPtwf+JyLf79bk6NeZNbGxzKiHuxsv3BULYQHkhlTqAkyZbxVKmkDq3nVb4
ExlDzJ6G4Fqu1P+DccZLnWMjFDBc56TEvqA9V5iWzxv7nCvYiS6bkr/2r1+1zdx0cseq5/Shxumi
R1KnAB8TZbVRY5Jwl2zPP4C2doad0e47fsbE3vdQRHNfRn8TD/FtvWP38jpzFsAgYZCfAlki03oP
1ycryrTVbPONr1qjNCmjDcpNbi2U82+Lbfr8wrAxMv6Uxrs9r7bMpJKBpv86MEDKsw+2iHpLd8Px
4OCKb9RanuaJcN3tKz+y2zT3iq5OuAGyyZErSJPuJBWn8cVEKv+J3wkkHBpfVt7GFSfNd1LZ3zHx
Z8qnhJI3CjN3K0dNgRcWAHX9lXj1ozRdKir3ti4eudGLXXwLgbfFwo1MTuYnVPdProsX/clJh6mU
xpNPjltAQkJ0IAFUO+mFThkUPviaGCyBlM82w3+IXrJhNZcBMFKPaXumwgjVpQN47h0aozkz3AQj
NGLdamxcOi13vTeFNRcr3W1ixa63ng7PMzdmvWXKMOrQAmekgLE8ql/hH/WfnbJ4qtQe9weUSYf2
a0U8Qf9waZFmnNyjjlW7ouDqBa/v8wEXJBOGhgNmQFv7kq6hiuWSuewaJRgbVJ+cCWV2q6KmrHHO
+kWBoBgRDCxV4I5N1THkCjO/fQ/FjEY/yrqoncnrbZNUuNyUYB88GxGIwccLLcSBXLCGKtXBxZ4M
OYHdBBv3Q5pFdtdPTgDwpuwhodMjyH7uADgWDlXcbmreZ0pNxUWaN1MV7bDRHt9uKA7NY0gVNJcT
46lDv9MiW7Ivfxv2o6rl/+bXtb+zSayL6mzhg1qnZdR8jgOCAokFy6HQCLxrJL28ac2MVftlchkH
lFB/3hlWyQdEMxy+y4Msx3Y0e7GWOmnG2JBM/An9RBqYiEn/l2rxc4YHondcJJFSZF/jXqVuq87U
9tmxKO4oEFx2+UgUE03rrf0ugrBnX8itvw+LGz33bun3xLVMXZktpmXbhrmeI3G0ovU+Nh40eTmx
g0MIdHb5zo3Y+qzeSNOtMcp3aOO0foNC4HF8T1byl5qof8ztQEeBrLGyTHTt80RwYgqYQtfA+5GU
lr1vCc8Zn7azN/JvGC7jYACMsncWXzNW0GOfDWpJBKZDeLKj7cSo9j2t19pjl1ximB7zRsXOUj0l
I9PWCto+QhYbV6QwvMgLuHaqLIYkXXleF7+iguBPVV9YHJbeFeW7FpUYb07o3v8Mzdlaj1IE5Z6P
M6ZLWSN2XE8DVQzVMJBB80orYPDIPrOMkbV1ECLC0wvzEy7AtUWq8/jV2+NgDB7FKXceoAOO9hCH
o8Mp6uBQXEKj4gB6EF2PcnfQjgRVJ4qZm1xyCr0FyCMXe6qbHSf8ZDJ9AOMJtQG0c2H2ZXHi6+zp
giVruN8BeEsFz8iYUZIfjRodgz3Oy+5AmqF+/q36q6qbi57N5ChtvRDVeBbjQTSe6x4hHWr1fk/E
q4+3GHMIXhMgKgJZWxFXPVpN3UZjs0n94nRTYBPeX9PwWEZitKSyA9q11gD5Ll4UXnUSMBaiFRaZ
3wCxlIGZifcHCe2h8GtKUcvLH8ds5ViLvEv/dAzpeYhqg+aa+fRKwRvMTDAoNzofL2vQUs9S0e1d
TA7YXT2fZOUsEpJUIwXVovf6xm50PYWUZsCThQhCDLd7aSOmc3p6gYH6xzDjELZ6Eb7vcnQtYNkZ
xmvKihaXkmt+d/yxLg7Mc/9YQYaWFv/gsKYolYyBITeD+f7OkvP8y4XwJvG0lVkOb3ZVs7e4I8Kj
z4V9NvKgW4nUC4bpwKoElkMCsS9jeVeKFhFSjMyvl04Y4WxLDqtJHnyuy58IbcIxh1zlOw9ZpPgL
0QPH4dwUuPfWVzDG9Rz9WXfWIAYwC26s/QtFptLAOKwP06TxCuwxotSH6xoCpH276IP58+RRXnJ1
0ppCM1eERUco03+1gmuJyvZCS7Duc2aoxgHI+QARioq2stOQ7HP1sSbcDtyEi31B+I8MnXG7QeMC
7+TnpyXaBvtDA3LSX0qqPD20I7qkB865EcfbLCMoKFkMQ5sWJ4jLgHNGp9e+yXPunXdHqPKrB/Sy
+nRg7WI5HS/ABlEYUwTCCpRYr0DgYOl/L6VWOGmcR5XXyF9Bcz91Cvpme9BAgh6LclYbu15BFZVK
qqaDLT8j+Xx7Tq7qe3bwlCGFCjTDzl7S0zyz9PX7mECKPi8n9qF44TfFhAOSGmT74b7Op78oVRWS
wy6PUbWvxg9REsh7SQFlfPBQnbqs64aF019HadrPSB9Hi/9gGek5kQNE9Y+FDePAbAehKyZUx+GD
Pg1YEn5TiE9NsRiaX7gD6Gsk9qg6d6AmpnVeeoj/nsyoNzH7N/eqtdlPhjT8M1EhKnGpfv/KbKku
kn19F19Mj4U8hto+FXXJouQpCHqYOhlX+PDx7MP8MyH1xubgldtIp/tTtn3lwsY81t78s1MG5BrB
nrG5xKXrH5KfXPo94y0QnAxJGrPlEFQyYwlqzFSeAMVSZQ8RFS3QPQgJVWsO5YmQdKzyiEbiM0Ev
vRrujGGiy43pWFgqxMI84EO+8dQqAq5/RCK6aKyzvTMY+nxchF/rjAi5A3yIkL+mdxrl0re1k9vP
UO6BEAYssTGVj3gRKzZtdE0edf6/HjCJL40FOyWHW4be6HsZoKMuGS7gMacNWv0uwA+b7EmsqzUP
fImu7dUyQWM/N85xO1KEi30gJjEo4ayGbdcLizdDaEmaC/zBl3nThFjKhvG/W9ibDfAWs9ixSjSf
jtcwQpKr9+49/9BCyxtcTZt4Tch+5fNaeT7/m8NE5Cbvys8IsUC5Hz9F9HPWcA8TB+JBVYTLxh0d
Yf/3JuKZ++NgavpCBmH+cPyq9V6fOZwwz7AMkIl1SmWFDMmCkUKrYzaLcg0p1/UKoLSuBB43wUlD
XRar4LKqjzggW0RIyygWKzdWpS14dArbOP2bBt6Zgwhc7xqs8yVYcTsX7AqNuhx9xA9Q/aNpPfQo
4DXsF3uodWaaBzLGZn3LcmqqnWEn2TlvMQN7PBKqLU/yCUd046so7RqMVa9yQ2ksPd5jdiUoWsBW
c0nKN0B10V2ca2QQf67DzBXiepMKh56xmWPhX2LzFVmM36PjAEdNE+ntfu+RBQ/nt3SNmBb6VpSN
3y5iSw/c5fhe/mZsbhk5UV3yWxtx5BtV9zy0IqrMWJ7dKbwYcvFL4Spzm7UNjd9+5gC0QLqPxWcx
5fP3jkuiF4oa9JJqHib0WAMs6v/2QmFJUnV/UPUCN/oWHPkdU7NEFEKqRHhqyICEgkhUCCWxt8zB
N8JiTJJZG4NLXMSvZiVtPjwLVKPYR/ALDs+/+9wWwbM3IN+3yVfnnfc5idgOZ6qpHA9FBLmZSCuU
wvI9M/m4qPM7gnvgj4J6u4YBpmgEtbYw3H+T/hyIx6culsuchQKN1LptilMfKQAAcGeMwUXlID5x
5P8bdb683ixTPuS5oas7bAEav8n/MRgL87/PxjRCwDZO4mnlcTsd1d+d2eUNSC7RTsy9kMTrCWIi
l5RptmOJG5QyDqIlH6MseMstZWwwLuka+zgqFRv5v453ce1TuRcolJQKfU1PwGyLv/KJ98GJXjd8
XI35qYFP/xZ08VFMwrcJoLpPVPX18BwYohMzL7glHxj+Q4Dv7G+9HrJr/GcFcpK+K41VsS2yTPWg
OvpZYathEQhlzbX/z5BM3ZWGkxihjPvHZQfXTvz4ZueKBvZZCsiHn5MybmT2inR8P8/Ffh71C3Vq
fCXUQMY8o6D2+e3Tf4UB0o5Ihol5+xHZoTVj3n/vT1bty7vjNdlMoYPhKhYyt8XpK9QtEnOz52WP
xjeH6H40i6kmqBy46K/arklocMO3ppGHagF9T8rdN1Spsegumqig1aFdQP93PSAaxOexlomqnac8
wCBy0C186hjvnRcR/kCxGhsgHyD4RO2vrTLyojqP+ECaHmHJz8Yl5y83CciVx6aIfb90zDCYd2q2
GfN1gdpJ+ifi8YH+NHTefbp2h1W6/WTunw0kvJ91SFfT5P/TIx2CfKWM6viUIJx2HIGBqA9AvFSl
a3wtzpLNin0s/1M47hizkxeMoBHQFuhZo1nWq75465gjxyfBoXjiqyeeq/8NnMI9t27k2YxorZD+
XB5CVrtbGsWBGlNjpRHck9TyGvHY8f1Bf61zxvhKEg+xdnvbLnDZuaEiPW3FG0+rWgtCPc9yE6oY
NkZ6zg/9QtVYaUVe7mC2C/6VJHGHqKsU0yCpEAJCVvE21nQpbVoFBZGkaVaQRp24cMn3684KK4Dw
7YRw/au5PMBH0ShK32YpFxIxbvQBzQEsyrtShqxmx3KEUnyUyqeMbYLy4HPvFHU/VP9TLNR+hE/t
Uw0SYXGO1S+j0waIPtnNd8mtjTVeT/BJkf6NGQvsbMv2dLVPxQ/CRBPGRvtXJix3fkA39pop9xhQ
hE5CucN3DEGiBb7+X3laN2w4MD/E/m5ezR/EUzr7B5mmVokMlTs5X18SwYbaNBtBFSXy01dMOqym
V0P2soLrSTU2YS8FBRVUv+iqdwnshlXFjWw8AsgIyv/fm2P+zA9CBYLDtc1DhOACoaNQnYCUh0AH
QOKS4HDpYoU80p7pQjWIONCwWENeAMkZ6gArb3F6tUKzZNIa3g6Axj78BrJVsDRoVQeQREnWib+u
JByk8ysJ4riLCCDm+VJDcX2rouueDh9AqZcaNpCFtCaAwcuN7JxSxRStsmhuK43PVRqBLLg642OY
QnbY+FagcrvM7ztlrXfpLNlC+oTToD7RGO7+aT8La14kaZa1p/Gx7PzjZppq221DjQF3kvlNq5P8
Zm4twJnfNh4gdOSOhbaygHH3uZc1EhMCrOdV9IyxXslPfK/Sg2HUpMfrACChenv0VVsLKFrZU7AI
N8T+kBs1BbTTXLw2r4TVrkcEk1kL6+bSSHgGXBL15nCCpxE1S+yqySmVkPD+4eOsAeTv8LnUgxOw
iX1G59h+tqxlwgnsrdWPGuCp/rEaF9pqtSoCXbkQUW0TwMNMZJKqMNFALfEDybTp7wkkCH1SgZ4F
pnNCbpWEePX3ZmNd4FDV7q6PHWxfNpE2Ut/WMz7fXmgEW//MZ4jAwoMOQGZyjeklIDkFU0t5DbOI
CxGvUOU5RaM/vufVak5xrKbdlfTxUAST6zGt54N5wInivFzZbUt+U0KXtkHUKSlBb08R2yhnGo9y
i6tV0FObacfZMPOwvH0XPJ0+0ZP6+GmPwk8kNWYmdFO/F9Rjd1DsSy2J2wnbGJw5KWZQVmva7o/R
hepJ7m7wXA4VBLA8JWqlIPGjwT2mu24m7XvHNe5vfrd9NkuT8oCHQ8zWv+rw4l/zyXkev4iBx9TU
CPsAvoHpuSA2AU24bpKsocBjMHhF3Z6zmQZTkMMgXavXSVpqS6x+wtSFrHp5I0c2YNzaiLGZfKym
CsOpXxgVh/WkwlpGknPM2nnEIKkJUaPK19sx2yufVXhufUzO01bFkvf+/DuA3A4l5ewJlKw7mpD5
B8V1rOR6qirlFHXn+lzaZTqCYYxhIndP4JEekHHoe36TgLz9XB5Swyw7yqrZyC1MK5CBMf7xbeFr
r+Kaf9M8a6VIF0Z49YExKctVq8iO9rppEBmtjRoKS6PYZ+CVorYAOZj1kJeZQamO5yWuIzAfB2hd
C1Ay/hABNiR2lRFNhJjRA8QR+x1+7Fwl7kmz/SwTPR/uLRyP3d3LvdLu8IOur5k3Q6Z0eRLFutdc
o3e6q/OzQHUDgtp3csXlE7B4OYM/yVIgaN1rsanS5xc7XFoNN+0Wrj7w6PycFyRf7LlyJSqCxGuX
eHMDbXkzXtMX5CHa7hmhiaF5lxw1l0+fdUL5ZE1tlpdMYQHO/mFeM0JPHOLhNRV9JxMgXayC9Vmr
oRzO5tqX5Y5YIpqraUiotg+914g/V1j0fw3r0fTL7bBO407oxp8em7A+red743eCI6APKdYd5q83
LcuPfHCOU1Ba5sVc66l8FL2LjO415nyPobrwyuZejJTOg3EUV8aDOQop7siFfGzSD/sN779WhiUs
mSxyU3GPq72BJCT+iv8EwFnmRhIdupevsWWKMsaSEzL2dTrEsDnZnJqXCfRM4p8pccuiCLxHSS5V
FZAX6WHRjrLFqqG5eUArYhjydHcSQKqpl6I7QaWRFLmgyl/SPpN812go1aEBzdDzah9J1talQGCi
I7uHP58kRmzmyd5f6FvLcEBLEDzsN2zG82xuyht2bl32BoBFJkd5fy4q6l70c821MIXhn7k102KP
oNgUTnpW4oQtCfqQgWKDzZoaTwYfZl5Kue86Ukj3ixtmu5qE/hKLLaWlL6fJf36/dfx1AhcfhDDS
CiO/nIq+4MKz8Uwx1ZB+joSEtxRXqV8f4VfDLrI3dm8jFl+x6Tl7nbAkqlH9y2TBZNV3hkLXMKYc
Ol8kFPj5xDnqHnZulkzeneE/ZNw4cwYRb7DmPql/8O+TkNVidvK4NG54usHCJ3KaqNaRim0eqs/s
YWdX7rOJ1urOVzWO/KGyi91pJFcbEGLByPwz5f0mVHsq+wkmFpz4WqjwOTnLZJXB7EOP0gC907g4
vnRFGLYMkJqyx1clQDbPpXkXmyMy/+o+1ORGJqoUzkmCUp7y3Iy2o4dMeHMVMULq94fnZbniUAxp
wOPJyJ3TJoieGh0MIVO/HUvPbczjRJhJ/AaOBO740dLbeq4Qnut7QamJjgcQ6Vrqz2IkTQ/bvZAW
6uy5152Dhl1X806oE52FEdsy0rs5GjCobmA8z/azbBXR2MbwfHFAEysoRg6vjCwXuHKvJoUI+saf
fRZh7LK33wscdRKFEgOrYsnu1gq2OVLJKgJHsgiqZKjybyjKVR5CagkD+ePbValM8yGhH4rBRB9t
LvDVkBUufmzCZWrkKh1GNccNQU/2RLWfey5l00Ji2igEX/nRTlbNvg+3SIuj8qDp8ERiLC5YwJ+T
j46ivuXQ764Q1i0s1lTo+5+QAwG606rmSjqxMmV7tJNhHYmXRKAti+vhMRnlJG2jhEPko8CgaxdS
L1H2zQGxyT0p6wTmGXKE9eyDJT11cdYlDeZgKDo/ZV0XORXkNqRaI0wXBkP1RR7QHDrAuHqgxdRq
D7LSfa6vDme0fK+uXzlps84Vjl5hs1dKK/weYdCJ885NpQR2QYRxIAextEEwcCJs/RlzNhXjeP4a
bh+d5c3vjR0SmdgZoSi7FuqRwBI7dHFXMlNujL5bP4s3xxQnbKuiiNVBVnvgPLhQ1saLm4Fpq1Mw
bxZ200/EWzXEZmK1VFo4eaXLcaNp9FOYVo+TrHD9CGozR2RB15rTQCm77R8SL7D4D3f88NkmjpSQ
eaywIKoSGQeKsVUH9cxXqN/zW8a5t/FWXw13GKEFsP/vAzcklk12sMUNx5YIIK2sqhXAnk6vonTO
LCGOBUvnQ3w1AITiWeaogi3YCkJRCMwjXBdEHgcgkqgwDdRrruh3GrVTsf1ye3kE4AgQXQjBa5zg
2jCcjUUx7T9LOTwOLPNB16F4bEzt3eDQcwFX9qC4qC9MKeED2iHhRoyom4iuASy+C0uElUaadpwc
jPnjbiIDbkFfK5r4rddQoeecKbSPrrtlKB6kZR+A4Aog9AOkAYvQ8cqkCQiwyZO3bWKkBetSH626
Vq9stK8PP5b+ZLK6d8k4+vo04lQdK7KOl4f5uOk+1ZRH5QEEJAMrgsLXwv68yV5HI7oawixNgsJU
ZPm5ezRLsYFIt42Hycqbwzz2WbPwRCrNTLuJfQRlOlHfk/1PgoXcNgAC0BFsF3kScgp2ixEE20CU
Jf+k0Q0WUe3836fFAaigTYsfSPluOet2I+CqtDZigPU58Iu/J+RuC442BiKxBqDVM3OY2hn/NvEP
zXVW2xJSY3lXJJce4eZcvwCHHjjxwkV3SLZQ+KkEHezM7xo/dFAQmKORlb0gM+zyJU2/pO4g+upD
Gw90R4dtcvVQZJcfTbJ/YL738gJJQ+fyJBytw2mVWkwzcq8C5HolPOt/ggsg1iU5fJP0KNdXrhhN
ER4wyYVIWTn1H2cigsClm9n9nVjblua2pA+8aovROCUYbIJHtORkUEVtwRAZiPphujZ4zts4k1Oo
GPjKBVwmn63uvV5FcQ6ow8awfJ3jm6p1As+S5bBxwaRZPuX/ywgr50OXxlHmJxwHy4F71IHKzPie
WwvBEEuCMoLH8QICf562CMW+MuMtgXW7u05X1QGqimc6Q7KD71UWeIU6au4LfVkSxeDBPxKcMAl5
WnLcudA/JfWea/AJjDyED26qWYscYf3xgmwLbAqXwVtbUv67w/6COjyH4PRlMxOBHzgVSBGQUquC
5rs4Lg1ZoJCXgI/+hVNLQ3ABGcPfYHrv23161QHwe7thH11mQoiBK3xJybuuy2baxNlgKF798ihv
LB1mlUeHD7kAXgVH4fdFJN/KYmvUPq6sMOufHrmWzz+QzTTIFkuA4gZHOxwFy1EJ7l/CcwDNRDUs
10UlE4XV87D/I/FqB05sDH20wDFR8USd9IbF0uFNvghzhy31gQg75SfylH0XgL8JeVSYQwTS/r+w
9GvSu11ZE9eetajHpq70d6O3uqWyzJzk3HmoNLrHnXZy82ZH0knoRB0GbWDx1X8LDXQJCLH57J0u
L/XHnm+t9mi9FjjK1b3CjjCOsTYWGegFOahQrIiFTePQ4CU4EM0Tj9sy2r7ZwNLwZBje6Ez7s66h
1j4ahdK1IAvWwFY+vzAcyEEVQ70v4TOvcawttq72G4XSn+V4H6Dsuc2diGY2jMCr1e7BOAafrq92
AR9ubUn1Fk4Q4aMFnJXMw8wngaR1MS+VdIAiBUuYQpG7WNITcPaP+nuT2KPb4BE+Gph4wb2Lgiw/
VgXhd8W5tCytZJnhofOr6tWPE6DAtZtllO6LSutcZ9+LLriseYc+9rGAgPO7B7Zm9Vj3CUMsJg3G
+MeTlB6mV56YEOR7yiMrjNcbQviQ4Mu9ZF9w4uXeaTANJ9TqF/IKJ6Xgr0MjgWyLM8VM/hmwpBvn
2DqUEDk2lnU0YSRn8QGawr/SDDGQg8wzqcfZb+XZI7dBv8swdhOaMIo8GcfGe2v8ZGE9j0HYrZEK
OfIQgk5SpUs15QGetbcsm+HIxyk/KnWtr7dA1b2Jqs58E+nBC133BNpkCtBsWnTN3O1RSXl7wL+X
KnmJ22UWrff4U17U8TyTuPQPmzzqbDSlR1/Wv6x3nZGErU41B64Gppy8oUmtWu+q52XHoB00lCPe
NI8mqR6EhgfYeK0TMtKOBRvk0uU2ISAG6SQBninpM1AILP0uGlBtUguJ2fDlZpeSzDZKtdqSBgHJ
MlKjHNeFYxH4VPq7QSLeH7EMLYWI6UGS6y2PKdSY7EcvoVz/9KJlN93PJKbVcLYJWaxkBmbFMCbJ
+fUUAD7g670zlgaRPj1OmfJIW9Cg2L/tt7AMp/v8V5EfFDq7dhjsaCevFvdh1/ftlMDJ2CnQIPJO
vIRnzR3FoCdiWtbMc2pkRl96dSJ5RQZP2NcPwyrRBca4eQix3cFgrEF6+bEqausfYIMwfqfJ1COV
tbeVKNyQORDNlFdPdqPl1eRWK9Tu8Hw9GPxZTsgGfy2RcGj50HiCdvT/gQ8FR3fgHzyZpTinxMxo
MVaaTHI+jBjdMVXD7jxq3ke/qT/tiLSkR9cDqow0JM1bTGIniTqJUd3Wffl7Ddl5cX5HN4uDuQ2P
3mANLe8nE/OBvLASg9QGIPR0mXSTyPgmct91bRHbif44ipzJiaZGCk1e4uS5ph9Iekvz0TrsO8au
Em6vKKcxL9ZKFkvx23VPU56crlbGgYbZ4Y+BbfHY33GJSs2z6LXtsdgx+3J+V7bid4MiviW9iMHg
Zm54f3LENtyIjxLYM6etgr0gHXKiUY/jLUq/uV/y4zfBmnTkJpGEC9Gwyjrli6hL7Qiq8+ANRfeg
9BgrvR8/jbaz8CW9ZdU0RrzSNmTzIkuUPEswg2Su/gnsbahGuLyOTal1vPQiW6GyauxBPxdHz3r4
wvn9pZskwoaAWH8eLie/k5qkaw7ZfWtrZh07CfjqepPLdJLfgnE2gAQQAgATxQpsnhnfYWQR2h3n
XcIeNi2i0wiTlrunnVR2YSFlW/mmT/Ayc3tY5/3iABDybQSbjcFlPn0ZwL9uMVyL3QLzu3JjVetd
SF02+iKEr+tX7Zt6X37+Cmpi0sJJCuNkpw8SomCjHaAHgL40xsOJXeMbRoMhhTcM4E9bcMdF3Axh
Vycouy+4f010cs+qlDL353f0ZAEMN3cQ82NUKl2WDgLQYqo7f8BTB2jGssP09lXqOMJaQanw6dxC
sJHJ5gPwwORg8uUgfozptoH5z6Iwv/5YDzH/OAzn1pbPKr7XuMr6/8iPxSaYgnE5Agg/ZtkOHAXR
G0/RPR7a44hzmQ5CB4DME/y7nJkOg6UJQJYqHRPxKWfvqyal1ghAur7olaghJQyiRi2u5sw/AwY7
jTN0i36UOLXPFaDDeLYkdJC1S6PIepK6MDjZjwHE0U1KCJcjgAUe7WSf7TSe87kYPKY4P5bgK5rj
S6BIzoczmF2n3NGx9o5IYGP4s1iAJglrVKGpX5JV3F+E/bD3JnwElKBCspPjTP7Yc85vCgJC5tyU
EooniiEz90F5w/+KnyaWYLaefo7sv3SWAbw51E0/VN1W9BoAcCQ3LfPtoofuBdeeHT1Ss16l6C5Q
NYcjSg3YaSGFgJbDasWTmfqiD/2DMhfuAJ6+O6NX8PmKGIOa4Dfzc/TdvQrvC2l/mUm6XHhWHmX8
x147uadN8CznGOxrRJ9r6WTZiKD604sRJwZA2R2nVCOpoRuF1HCltL2VYWi67J7UuEZw1qAJT6Zu
Bn015+at0c5+FGWkmuwmB1JFZdRd+LaHx+w+vsbGUm17E1Uyim8G64lsrinhJwoVfyWqSdwx/00C
lxNGBdAx0RIzR1owc68AVwyW1OV0Qg+n72uxJwJYJMe/I+nSrImW/rbnzHvwNbxMJuI/qF0aP5A6
SW6rzYYk2Go/BmWCj5C/fdOYGb0n7rsn0pTWXcaWTJE1Pniv+WXLTZpDPHYPqQyq6IuEBsY9unBW
zUmLGRVputy7/v8OXfZVnOkIyGaIsAkRd7IJgIiwIGcLQ9oD/pAXMAhBJZUWblQdcmasVpH5PIhL
sA5C2iEn6ieHaWbduPz4LkZFYokCHJqStVgbfN2ZmGrCuIr2HA8NGcFjt54XbP8yMnS9D+7eieWc
ONzkXYOOFazvNrR8LIlnQjD1bfO7rIzWN5Q9hUf8ORoMav3/G44w/rdr0OnyuMb9ioUapTPmrPyn
KbM7cS9VNyk4Ik241nCKs3Y6z4S3HC1ZYcnxtyoeudJt+45lVlUNl7NecSg4C+Ho1mpeO8AOzhQq
Dd5LSuvmcSro3O/yB8PZu5SzvmDfzSPRLM5yJySgTKKHiWkmrhEvnChbyaONVGB3B76G2DiEXsuZ
DEpuy5auvntto8pv0bzarXHKNEM1Ft/1q6vDmoT/4hF7ARL9hhC1tK+7dqpj4HwU/pJ7zBJFZY3G
01Bdm0xcbcSRbWAnPRwLGIk+gg9lMvBcubDI3BkynLVgFROkOW7S9rhj5R1bH12Y7i7Kw0w6NgDQ
Wj6C3xbONrdn8BO/GZIjwrlN8x/BGdF383w3kpGGhscTmkyhrVoi+Zd9G7e9tdl6SWgKLOX9S6Kj
OyhafGB+NxStcJRlvETyGo73im67CCod9TCE8aQPzZ38++ERAi+9Z5kYcpfFpOyu7oX1HCYpxy8g
1c1e8mky8/Ez/oO84OYQQyZDgbV+BGSAgEJknw1oQ+6OeX3su7MNCGYHs5A7bEGLyKDRgUns7dnz
y92ICgQyzPcrWMTGIBqqIS6IJM8MsF3rAoqX69aBicrZlSOrTuw+v89j3e1wleG/VJhBxPY0U6Ib
qeYtVKDBrwZx4Jf5NIlAdBUVH5oPLZx4iQp8v7YozOpm5NizRfNl/Rjsw2rxOWTIEquL2yMmgcrw
RCml5vEY/IgpFBuXp+g2od0oJADtL3zckekHukguGE4UfE1X+lDQViMvNyu5ScPp30Mj/5qIqT5d
rr2hDRl/cLiw2MgH+wCUJnBbyCMjwKNoOjhcbbNNQTm/XUrfJ+XzMBVoQktMVhHv1COcLJ/ftRMA
iZCWhTs9tskxdlly4fDl+5s4tm9PVYzomSzlvb4lt76elbvvvOXVqxCEgNfRLVmrWyuZ+goRY7Af
IH2HRX56BzuqMb9Bm96iOASElkzpQVvNl8J2MQZlcsags9zS3jzKlK2zZLAJlhYRKpcEaKHog7ww
DhFoxxMW76upO6sgqxxA3LAOGhPQGqDvEFrVnQlEUIiG5E1s3g3ft+9FZmnW7RC7OIK9kzXucrr+
0qR7UO+7SE39HeXWVj5GvtDH7zrwi6KmkkNUvrkvlYqAal/jN4HqebMAJR8GtbIDllTwvKadXaTC
8m1YFGV24kfS5yVacyKI33iXUWM97FmDQhSL9BHyH/kXwQtIerF66vEDmkawqzvbtFIbxU9cGzMl
rY1tr7EBSKi2Wzm/CEAquJI9xMLqx0dVpruPvqMcscasDdK17tBkwQ2Cy17yp09wSsFk9RG/XUBt
D9BR3fWtAF3otpcQ+s9nJAiCwXku5Y325Sj+/JBAKNJ1qQulm2khefyXc0VkgwhyjlmB16OiiNb+
w0abQYF6eEoVe44H5M0go9GXL/dxKT5dmUoBikLe5khM0WdMVQeOaailEh5siT/9IJLAeqIR4puR
lPq+yA1pzm/s26Jb4+ZRyAl2rGAI2nAEFYX/WoVlR3rQeJtV6g9jCO5SBWHGw5EqEMVPuwkWMC9e
lZ9f9YrCzFOY0Xr1HVzzYGTgxcQNaIeEh+GLolTSXNcu2xa8+gPn4Rpla1v+TZGlz39M0xMYm2Uh
7YaKXh5WG8ql+bsBzUxsS+UgLcYKoqCbc0Bp6Rf3TPX8F0WzMJ77MZG5TbOjLOEdChUz9hvtGETT
2rJtaJVBkOMv9wm7oz4ve6NYhmyHnndziRvWNokTUF9Cu0surY1IU3+YfmrrrGhbzBqh+/oemWcU
nDUNaDFmcN3uB0GFlv7Wt+cU9OhyzJ4QdX9YLkqaLy2aDaD7JX45j8BCwxs6DzADvqh5nzoIvvVA
XkEkc+PvzCHQKlBILJPhF2pklzx6mEhI1U2gKYUuFljgOhZm6+p7AWhhXbzhFfD8TyUXIVbwvurG
5En8ArdkeTBJ0d7VGxctTYBEvGBWOEcNs7hKluePPXdQG207Mr3s1sD23k3Mvq9nzg+EQRfnxRrY
XkzR8keCK9UNqJDTu/Q1l+q0Ie7OjcDnu3QsMUau01VjAFO9TINK2rjHOd0BRU2pc5ClT65lpYD6
2kqos+l8+FjsFoGBMm8ZLYhORew7sCxZBV+Ue+RtSsOKPljg2V/Yv418hea+0e/eZeHsh4yhgrL+
4Y7zQp9zHlTT1ejBHuXPpAs94ihRgjopPDxIhkAaGYLsZG/6fz+fFIf2rDQ3Nq64SWYfm8RqTFFf
ju/J/qXh6TtHWoNbxR/NCe/Qtx7sckJ1OhFAr43GwekvZ5TXdOVTAu+QSD5d9MNkV7KlKf86szLN
EkjRZhpOS3MOqs6Sog4hO9kCgN191gkaMLFo8bzy7SLp9WpefTGa4rAiL3d50+vEde1SeBUgPiaB
gVuQWKZNyd6uBV4tRPU1Xo5CXLwrP5MTlDdt6h/yH5ayZfLLmAk+LzVynNTZm+IXjA2zkAilloYk
FKgq2uC5D6DQYVpaxtXr7OIYSSKMK2K6Xep5A1VAG39I1v4EnurdMfmAVTC90RTjek/HRXueA8Am
o+43sT2pKI0Xmkim2DiIDJS8A9Bw50Z6VnZtTQP8Tjps+uPJG4+2LzIL+BXLvxdRCMsavofShiBL
2/jTYTNrb4+TRrBW2RgONFAZXQum2OUaII6nq92d/gWSz5OWVgtdOdCm2PAXC+PUrp/QU3rcXNrL
0yJEunnuTtT56/AxgnjAMmU0FW3ACtvc2qzSw+0m9GUgQVIMdcxcTZkczvTeyQsKqA7lTAGnKRNb
vzhgpsnqDm4Qq7JRo2e5o0J3lZAEzdQ6yzFIR1JR13D0fUTxt1bEs4rAsLY7NwyC9G8gCfE6w2mg
Xbwoheru719n0HtR9nSD/e6WmOANewz3mX/LliGnnIzh+wJ4wDcZwtNe9L5n9ABTx6OQgt6EW5Ye
d1moG4LG+xXvAi/Bm25S1dXMT5vKn7cbWtXNuElyzIwZqoGilt20dRnUIYy/XAOfA8Hwzho+HAyL
tzy5aVovvaXCeQKcpUWPmX2QHyha0sZ1v6ETzocafLt7P8kvdUI4ijdaiyw+QhftTuoiVIAKBPEP
uXAnT5Uv2No8ye2jdHGYa3lCtuR03+hwrhwwUohVWdkyGEHFEj+H2ZPQVtcN5dMhBTD1bmyE82OS
6tFLyzj8RVHQT8InkqOGxa6KSjdxQDa0gG8awMCOhv4m88U7t9mghNtLajSxWGb+t/zLgjdjMtKQ
XSjIRXFo5IaOOGToGZ3DQTzr1a6b0qI35U4AkbWBNmevNMZia64hQr9dalCwrwnfJOzIhXjlJcow
EQvbiPWIB66G6OXpVN3XB7a8u/r4n2beSzTpYbbmICghbtVret3Wgn+Z5/BqLgWAXJur8S9vkAtv
BEW0UV13IodpS3/kJ1uSTup7DSZFtgnqKYbRdXKcgu/6DMSeAjB2urTXbAZCuovnzonPSvMhoi//
mEJljA2uOGELlm7GuyCr4f6YG9ojZWMKzYeqTugSIwa7gxB9K8qIIWnsZJZ3GsS5q/Wl5xOEoHGI
zMP1Y5WJZ3/QJGrnGPoiNtNf7i95/xnE1JbG0JqAoDvPNYk11D/e1Lny8dqhLX+Z0vWiqOYIq/Ky
qZzpP2WMh/C4JJQfN4IhhDrUva4kvXd72IPiUsy0wE/U2dmYa3Wz3SRgb+JA/MsF0lgmW56XcBW2
MwoDr25xS41ZM1llGAavHSh83gtOtAnytD3EDGpcD0r/3NOyt1bOhMTipY3SN4hoth3OLi8H4vTR
NaWN6Jg3hjKpaxYFIKHPl53yzvjuW+JgDPnq4pr8Y9FImW4wxzjTH8tv2L6sKK6Nm4WlgwysAKm4
+6SdMCLfQmicIGJTSTRLrFaPtkWJYiCZlChKTXQdeHmLKvS25ktsCQvSoLKxPCT7JzWl6eICOkZJ
G75evFB3wYMrEBUxxI5T/Qq1kPh+PgdND4XdAtkAm3fImbVjx8KnwF94RjjIONg2p7rW10TZp5b0
VILXOkLyTVigI6ZwM/WE2GoMuuhBvqAfuQoq6/CE+x3X28d6m3vnXMAKII19wnh5/7GAnW9ntPF2
u5rv1oxXiItdXFXMTnj8HllPdbANlRH3mYQvBidpHgiv/7pvTFzr4Tb//EEkVtICIviSQNxFi7Y3
FtTNdjTgRjPkyW9Acja3nvzRwxIJOkZnS5RMga7WJEVdnJI/abQq8xvGG+RHRAcw/9HAEbsm7o8u
MuF2wDHRqV6gM1oohaj0OfEHQ2gfTzTjsCpjnIobGjawZ+7p/lAHegwBj5HHONrjpxxYwdmQPDd2
Bl/fvR4BL4KB0ulHU+E1AxSqK8lJHAnP2UAaEJfq4/9Uz3c2CTSHU3c/haKftKPn3/u3cZ21Wdjd
YhilrcCbtQZ6LKsJsU/erzWH0wa+NoNV+81l/KFJdu5X5JvWWv0Hyk0tpsHbcTS6X5UmDMGMNG9L
G9RzgdaK0GkyGCIGIMjeLPYRJRFVCsBhKQ8MEMJI97KaMGrp4K6DJSZuJ0Qi/Uz2XzRROe0bOUog
C4rKN56XAKWqxT6/syBhHOhGfxvCrIsU49S7uM8aGL+jyYp5BoBamaTL/JhPJdxcFPQdtB42zrj3
oAwO3KP3Hw6bhZuPZ++zJVRJDRV3PRosU4WlW8/0/vI1eZ8Hy06NPXFFLHdYlQMwZHev5/EA+BtG
DKOyU4KFAu7Yda6YIAqaYxPUqNJEocdSMVUclvv2o65nF9HiY53gLETY+Bucl9captj7n2XtKbNo
kUe4qWnm+1YnRjoUzPxuYpL+b/PwrTGWKeED7femG8ry5F+Khqjo9LE/4D3ZEWfnmDaz5hxO8vkE
hmzARqYoCa8smpKerV+qra8dmP8hwlsSLhG0as/Ik9JuQuGYpcXZv0Htys07pepXOhYCxjQ4LY4w
g6Q9j0hCsFKnIs4hvjyDEk9tRsmMpslwNX5R3Qe1eiR01etx2C31O3NlXk4maB2jf4SzGcHAdjRf
vnDJKO+roNMJMKevL/tfQxAdw2oF3euxQslREMSvLy1pLy2r2Pi4ljbdGmY4kxnszSxC9chGBiLV
QzqjecjKj3I2JXewiazE5HHsm1FCiuxI4YycM3KSjWfr3yonQRFyVGYheNAKG4qx7XUbyIga6fl1
1KaJ2uKHkOQp64lfm6nLna6bAhSQlt+Y60abU5PR2n2LiNmCBwVDtSZxnJREKUU7dCHSW9KuSggt
/2ds8QMKvQ7597QOV9oNhjoE5UxP80C5ieh2lAtJZRuHOJWPn7IoROlnrbLhX87YxP0z5AJG0uKQ
H9RiJKxI3mfDE7MCfqYmecK6ROv/6HfIwFZarFmIz513Ez3P2Nb+YVek7VbErJKDkfGO74jXthPN
2Dv4l8xk835VIbhx6HtB/Bdr2TMZar+ECnall6umHY/ou6IaRKYuqD6a+cjrwZLH+8aD1estUfdk
qB4VZYd/XeCnuQILrbEVHsgjVbWelYEMGp8meijDpB0i0j3UFghxhv02r7itB3A7S/PTBHcFYQv6
b2ewrwyEYoARi7z6J/nDtSv/p1IHtWp0a/0/hrrdEnTBUy/sGjzdFSza0TA9u1QetRvlpqQ9Hl8u
lFxkQo+e5W4Lle+STvmP95OLI0ho7E/CM9p3R726Ylny+wQRN+90580TPFZwfzfUvdX0Ak9t5ELF
7WpcobAFCSr9cawapqJqT2fsZznphTwyw2HZwoS28WITvkB+iwfWEPa+GMEkFzmNuim0LXBxf79b
DAmUhJrIC8zcepdHspJiOkefWSASEgqAvLo09WKQDkoo2tac9bul3Ir2SQElWwx+AsjGoCQjEFyi
YUUsy3QU4m+rrzVgnEHPF7Ae76Cv1c2pzVJl20OJXPbqIbOe6HuU8u5hrsILTG+cK64glTXCrhGC
DnGtjZxhwjFXDQpdzoPkDeuy7Au04bnQKnlEdqpYjbkOgrEnx9I4CRxHWpbmwbZSxos9o/pbiQ/T
xD0Ali3Q8L9vHqFeUVu34Y20thsASc+m4gTfB9ihWfvn/3tynnp+QzOLTPQB7+s70scGHaSK/SQv
j3YgKpBP+tUgfCvKooXXXKHdb+o39HmCs7xpM98UNivMI0dTRhmsqEzBK9F/WaYK5fJamGWrOfPQ
2TYDZXWD3Zz1tmmr/LecxBHoM0wUk5psKpvyxe53sKdyMEUqQQ5J5U1ddkR/cMjUGqsuLmtyBMpo
YSGgOyJ8JUjIhbHLaW3hgjk8bSftqbnepCbfG5AGp4ZQ5Em5dvxp0i3pOliQM4evAFJjH+YZ8u1U
YrILSokOfZxAMFRZkkp/i3KbYbr5IGbjx8nWXE3b9NA6XW6YnojGM759I93rQTOS+E55/kmtk72f
xDJJ47x3Fgl9MOfstunLm3u9Kq9SuODLb0RCic52Ig7RWS83mBA0GYZNQTEf1Bk24gMcuMyo6j1/
aMltNBG1Hv+ob/pxhSLEDxVCQif08I1A6U79UfURc80a402kqeSMW6EMqm4zBXYWfEr2D790muve
f1vBKRw1Ztxi4j5+jk89OrBfqHjQzyirw/ceTHx69p7bgaPxwzYPzr7Fe1HR2eSXyADdiHOYbTq4
iYx31sOVCnEy0qK2GBvrAdbaj89Kra62HKFQKAJ6XdvpVu3LOAT/PnyWNHrpaMYKwMTEH6V2T76B
FeRWNxaE/oRrGJsWyX9uDQ+lSiuG+nv7uRi09TGhJtO4xcMVazIW5M0r+wxNpXznbuwBpA+sPrAj
+pRVStoP5Iis5+7jiK7jtkxqYOY2jsIPACBzvKkLc8KN889hYy5Zy9cEiUkH2K18j2RkexejxQMY
IEMimsMO37sb1zGbJSIRQ8fPXXX1glKJ9RTVeJQOOnYQwNJVXpuGOrurFp/T56E5bibJNtLYYhBf
MOPsOWw7dtX8swzwo5nQzb5J3a+t2w0yHdQGB76Sy5BENdYLGl+eTJNo7BrgpAl+kSnkxcy6u49D
2v9yErZncozRX+81cWEVAaSY6FN0nZMPLmHr+SKNdhSPJ0KlvdakjnTdOuNXsYzockrZ7b9/+ZMM
EVx4UaqiM3xL3qpPKIAnBsEU8sCivRIVsIoYKLSDttKV4HYVF2cd9eIuToTaRb5TSsuAf3G9haRl
FUiV/OxHwpNT4WO6MiuuineFYAL3fJdWbkzZnXvAuxS/O6xT8tMxPvZ4mX+oHmS0j0hgwA1teGaU
v3tJigoHrbiPIgRBQmhdrgIxeRBgqpRYu5egTS5DHYiwqDMf0nV6lp+iXXTQHycT3n0YvgdFRIVz
kuFBemhN2cD+DxmXbwWHNmeH7wcRKXObPrKHUkECpA6w0RWHO81hnzQk+DrCz1PtF4ZYzAcabMJ3
iadNmUoCGI9jD31bLR1Qx/yuiBVTfhSsJUx+UE+sJVLLaXbYOf0D58kQS1ob8doLRK28/s6PFNhs
RXH2CEcb/oFmyXQNOsw1CfFr2ufPkWbW03I/IYdkszzxKRhRUHHANjuPmmrreIn7FsxZs1qhEkDq
iuXqdSlRaQEk54XYDiCgaA9QajpWIgrHn5iqgtJd9J+XzF98IPOC+II3UKZYBNgWWPERqyik+dD/
p7V5vHnzzZdIM28oBdRPu3y4xSjv4Q01hWl/m2JXJrHTrJ8AguyTR+ZaUAyr76PDlIp9yAdzbwNJ
UFGRs7h/IYTQQJKXueK55Djqx6OLjnd8Zx+9gfQbFkHnkyzNkFNJF9fmPN+36ES2QTQWfNF+8ese
4mRDg7EMzsnan9w0pF/NQm0AKO1gefAG8nWHxv9R62cm2R9yDejLj47eZ+PI4Y6hEV9zviZ+i23p
Vo88GKhI75U5QRWg1hYG+JNmuD4Uzq2uAHrVKtpg3lnwZ20JVZp7KpR00gohn+khsT1PGnLbV7Q3
H1uMoHVux9xCqzoT6FB1jkmyu6qaKpnT5TnaqSc49Lx4tOL45Qm89+Iq89VfhgLXxuviqCn+QHc5
YWwqu30t6fModdPzcNkUgo3XF2u9ehA70OBvnHJfEWbBmbMknOluV47EnD8PCf6u73iK1CX1uRYF
QlvPFJD2R6N5kP02lMEbCYaudEj7TXFdZMS0Er1fzlH4nyN9Vem7FvmGTs+2XyaF2w1xAKIC85Ls
iooUX1T/MOv37/RyiaNyrl2gMd8pxVJ/a12h2PONFHhbg4V1DAI13UddV2E5c9h9icV4IsE1TXYL
h9clK1c1+i9DBlOUkFTyDwM9qXKN8PBSh1GLdCTkn3k4sDX7E4Mb3pwrfXieCvAJz0rmlEpc2pi4
+ujGjphzHg9ctzEVCmhkM1adrCgZEgXTJdRTFOYxtusmPvAp/dU1NLXzD13/Hk65qoaH1yh9bQhS
kExvts8eoTwm4KCFFmlJzq+GOviUYNQqFCoHJgKWfOhm5dV67TaRNklElSB9QX37LgyOlM1eyzjx
qDEQ05c7I+PJDnsYTEUv5+JwFLqrrFPah9CjLoOGnl5Zdk9YQ5YfPZRChAbq05duQMY6yzEe5tKt
26yecyc/MOt3y+lGqQWVODkgxCKRHyQQHFM2M42Elkl5DV2pOrWTOazFrrFYchtH/CX0LSa1GiXY
Nkd6ww+6aUCQIt+CIRi0RmloPrvLLcZwWkas4cJHwf5MBc1LcR/njMuAppA+teiw+CsyVmErMA7z
jtScHlxKSEJfNmE535RAB9aX0qmyKLfVX/+YqwZ2bmbiE/ZoynFYGomxmawAE1sX8DuPF8gVlXSw
Zyu9C7FPuVm+w4rFHJdc0oA7nGXqK8Bkm/upsAw6OkNQGHtwX41y4oQTVyDQGJvR5yIfVw0JB0C0
jcTElNX7ZAr5AYjyDXn/nwBtqcbTYtfjEZQ9RMaHlHenkKiBdlYFGrpW63dV2OGaDr/BGXYaELxn
StMufQOcRVz+2nulcxtPQiRISPg6sLs4299r99SE9k9n51jtG6Ttt3fzdyypBxzsfBLqjbnnXxyD
4QeIkp9f8/CvcwID25F+UuwuRghBewC8ujazWnwGUzG5qH5+XOeGu7uEHV05YY7vrQCGw/pabHlu
FUok8KZdxqbHfu2eaEAW7wRzntm1otW6X4u0A1BfrUhnuPC7ZRezZETBVfKTSt9JDjZ4V4Hl3lex
zdGm/0hUe+WBW5vFoMi5PtmcvGERB8YAKYG126m/Iuk9gAXnEJ+UrThy0R2+yONlhD7bpjrqwuvJ
lVXERP4+lf+VFiRYxrl3aN2N+e2wunO4KsJKTK1S1hhftbxGwfvqf6tuLY1Up2Yd87ihoWLATxVC
a1/Fd9w06oxykSgp30rNW4DkT77MKqOs8YSE4u89/cjJzHxK2W3GrjSrhXYexCV+ZiBDpM7wgt3L
AG82My9GgdsXaWqQOv+Jaa8gp0UhLEGd6mWf9bAyfQ7rpsEltdoIA9rh4TPnADDEVHXfODa+/lOn
6/m3S+M6EQZgfWnX1wx+D2r31QSIhSZ/ntJttL+WD2YEET07RH8JQgb0/4H7qLBg9K6rnAmhaUSb
8GxoKztl2zYWJbkcR8u3/u6eYarTH8A5dlA2vR5azbe2n//1N6Jx0Z9QFIUDI8YuwojSNPspZU7v
8/8G7XVNqeAcI2jNdxFAOxYDQGiKuA/7RIXGzdE3/bkwsnBUzPpWJ5zIwZquNjz0GbpJyVOm1m9n
sOKY1/DMcAeqi5/31AeEb2P80GtTX5f6jav8Eh9Ul+nV7BP28m1bOh5j1KSepwxo79+P3PCq/NM6
Rvs7l0rlmtVTwxbapvlzR0A89XEr531g/lsNzlFwn4Q8Q4QuA8hia7Blh0cjb80o/BGO2E9geK8j
Zs+HXv9Th9QO9Tk/FI0ojHZNYLEDJC0J4H7Ozddcjm7mMACKqgHto2rlxFomMM8SmDhpsErueW8Z
cegXbVG1U/u2BODG4zOqx/aG7hSWFnJTzpKzEpFV8LzINjZxXtF6nSVcp0Ridyj3ve+p/n9YM+vh
grr9i2KhMMyOhV5PRz5JYVN7xiL55TmOLsikRyHO4qSZqnG0ZZKRJ3//6WBmx1+0TZRc1+VAafeo
MNtj24YFaM3lRnvDbfAtpdtcQTim3PlPAGvBNkubzhb1OBnSPn8AXQeJdsUJiHejq00LunfG9D1Q
y0cVM82OX4fzDlg95vu8Ye197b3nJAofmLkBI5AVf9Q6elC7rNO/S/RQd4EacWZI83WXSfSsY+Po
Io21IxtR4D11cHUAIgo+NOSW0tfg28HrP94l6doe/I3HhXAtnfxBuX85AB9jiwm8FjQOyHKb+0vm
6npVSwVGsXu0RIzk3co5QVzYIi3rCrtXUrDq0opUE496ciPZiNvI9W2v1G1iSaHTHVg/8gVCLM8Y
Zj1CVhcKz9bFhKShlvyjmQhbiVf4yu/mPOV/5+7peKqPSthMm5hxMxdu2CvwxkkLf8Kc3lzPpIpw
wdfAMXgxiw2LzrcAKKeWx9nNUvYi10iJbS14/ALMXZ0pnQ7vewIQS1mOyPDv8Cwp/hee8qgIsO6p
XrZBv+/WarM6iXc0evmyOFhQ7nkG8hqzyDIe14qXimmhF33A/CKsberQh/6oaTvhu5KZVVaqh2Wf
5APgsr6PyryHXh07o4vmELx8mUpmmeMk2hZDew4SXTD5JGkCSbuB5G1tKbW4djPjeadoWMhIRUc4
ASz/GFNU2a2rF6+VUY/XRhxrIoBkdWKWBcy8aQqJMDJZCmvVGol2Bc9yi2eCb2INzMd1MRxaXpbA
29+CijWPDbr9Jj64WswcobLPddfOayYRD6WwNUoyoaPkTZqZalAF58cLbI2gokGWVDfbqEpN3e1B
2nBoQm5Y1/xHLa5JJk0u4BaU66YEmWgqyu24vgONNqauEVMTRj5HktKl62LawpKXW8JT90TMDAx+
YngZRiFpoGQV3axMJAM0BBFGESy1D+k9GDm3D0zDCuvyz5r3z1tbtn4/9+IF2ImOcBHx1iOXt1+C
rVEBpLtg6fJ5A+Y+ovN4UkGIX6EX2XH28zTAIoe+jXe/ZtVkx2cPbvQPSf2mYaw2+SkAsoqhA/Ao
qFoWYpsYKdZhvpyJwER7yR3xs6QhE/pGALdBhaQw6WBjVG2Gy4/hl/WbNqTcvqHqtV6nROuKGxZd
F3K0OoAQSONawG6ScyHtBLcTNaCnaDiZbHHX12A3IlMJkWMjcLAvRp+Zb4eFatjpgRBpCDnck8Ed
bXQQw2Qgcx0s/06keAxIyvBKC4q/0ABlKqlJgtFODNdN73hrXpclz8VkRJ6sKkNyZAx5abnY7RWk
kjOy6Zh4xV3yw/e2NqnEiyjH7u1M3XqgrFVvyi1YKDTNdST9/yJoIPVPsVhcQuytydberjrXSJML
F38iYQkBsgwcWZfhqPkuKZRulgh+IqktSNB8f1/60Yktr3UQSlaU/LnNto0RW70E/YBHMDJCA5u9
5HdvSthP8ZGxuqYjXo/Y8H22vWZa99RSJD0nYBoWJgUHEz8QfW+3eB2KVmutseRf1l0lZc61ipah
dWw+uVsDlhnMR3WHMpWlVA92Kq9bB90anCz4KjCDSOn3bzxRc+oSRnDnc1Mff9Yo3ZjZsDMHTDgg
Z6snHyNVpVHk+to9SVXnFiN716nHx4j8AglNCwpz4aXktyRLhRupeZpNCfoT2CQFxinnyDjx/X7Y
QTTZG+dAID9ZN+SRtBN8DQCK8qtPWn9aVzoiXJ3hRr8lh7aFfjUIBuxF//ACnQXjWv91gnxQYJjW
NPVGrHKhz8ocQ1Pje5WCPqizCEqh8XFHY+uj9p75nlClph7GNWlapw8oeivkOut6PiRDvwiP1uAW
Si+L2zal3ljb2X0lMm9q9+N6zyMgiGVZJUhl9JjHlyE76OcaP96cGiEZlpatxfD5qtgT+6Frx4IX
C3Nuou//dTTVjvmFGS7AvWntpt8XDJ1ev9yvOl9SXY/uLgW+JnyX6Xei4+/iRU5MORH8pONcKiBR
obaj2zQJEKpJmB+x6WPfLmT/0ErG1k8aL/fpCD2slqCrn8BdFu95gNdE1OVIUlhIijeE64476k4H
R2ZnJAO+GSu2ObELi+Jrh5WN1bHCxFBazGUjUSCMPdb+vp26PuULAQwbt0f+K02xHhYh8e6eNPx5
8hvd/Pmb8BTzNWbDgxk6zqalgrva7Z0CuYKaVhDAldHNnmJoiq2W7pJKjMIun6WcD/fevO675EBd
AArygzyLXYScvGsYGyiTVthyXFRdZaHH8OtCMkYfTYXUk1mNTCgThyDh3CDX3PghCURTKlRZ1m1r
i3ZFf4xeUAqlEqOqg1T2FJfNofwinkQ5wq3x2i/s1dDMAAD1OZGT9fgOHZ86A74q5/R7G1/AxGMO
0CEsGIbm44lFP8ABm+qsuGKX/4CiuuYijCT3vTaSXh2SgO4+u2IJdhm4AJT6zVKS+ReeVlldL7XX
IlEjGtnSC7EGa8BHiZW5LmvAufMJUEJW/SWwssoBsIw989eMMC48p3VJ3izhyR97ZF0LXSzIL563
n6r8Ta87ZL+eO/QQGQ9ToLxwKqWyNZdg8B8C3cbdf2B8j1N21PX8h683a9oRF0iOFbChSD+5NfuU
exR9vaIxPmRLnI4ERbpQYBnrTna/clmLu7Blz8khoZy/m03i8A7a3yQLCVcXStECSSI6eocs8m9T
cf3iNpxlgCKBvmhtBx+pC5hi6VFnbLUnV/OM+oSa7uDAt4xuRMDvUd+dNnfJyII8rPkYn+ZBzM84
ylSYJ6gMXZ8FnVPfX8s9zhyqmQUJbo3NvaIIntXdclFlvAGNQwkR+2Y/GRgbZpt1LYUyLncmgt80
ZyjkMKxqW/oAO8iePrtj1IQ+H7lzV00uZlqdC2cccxDf+oOqfw9XpFxMrs1eWg+WWJWPy/LXfxLX
MRiiLJo2HvmsAZyp+9cRfhRt2IeleIMtl5629ZOlYFWmpSsIf1Z6LeU9eSEXE8d2TADZ50KuybRU
D5i5g6Dsq1U0vA+sgX7yxZI/cSdGzhe3WHoIh9XyimzgPlP5Lt1H2CuFb5Skp3ZrM9TVYBSYJn5C
/dlFEk2VtgOLrIjmvXtK8ysCpI7sjhU2iJ6PGuQl95HEORgw3pvw6DcMNf+M/vPs0GqnTbXvgHfF
DNZApdf48su9jIAHtyTrKwRWG2Omg+z4VuR8LxV6PL/jrw1S6FtKFFVqd3Jj+GzhZ8muwsxt4Mbn
6vl4MRGqlCtlBpDlZpxWonJTCSmk1bYWnLOq2lf/jUtvGtzK2I+oH2AqhyrjbP5lZR625mIEz7JH
3kXsNQkk7vXNzZfbLFChO3LFSlGfKMHBliEp1WOiIWmxr0b/Nx6T+g2u8oDI7/KK9fsYt7k6m35k
A8EhkulKYsh5bMGSdSV59viSzbR9qRl/J+/N8X/S1brf7Gr+MLhugPvpAjTh0nzw/TZomBSQXec3
k51UXHQ2FDWCAMhs1uoaYVsu3Qj/N4AC1cM3nZFGH6HYAdtEDPXsBLPcrV42kbGrnC6lZceIRmDV
qOqr1ziuDEd+oryz/ncRtAc4n8xcM8QDCkqsw/XeH3KJ9bhFkjpprkMt/ZqwRW6L5Ua66OMOsiP+
fU+6qFdAdHBEVoBF9mYEyuHGkHCcRZFheRaLQ5LeepnbGGVnDYHq0etHmbhLeqBLm0AqxiLWegTG
VR2Re1SBhu+OAYEFZ05yoAPJ7KE2449nwvM+yl2HnqHCYaXp6h/rA4py9FroQWGo+rf0HRyZtLMb
zb4sO5cVoNULxhAqAbCN5sLqc7LT3FGBxXtK8/f3+wFZy0lDOt157UMjfDxgYkxsACtZwUcxnAxY
zb+IkwcqWIQxxLiln247na1MO2aV11/ZCKDQolbFq4oHZgRvmJFNi6uQAF5T93n/CRFjMC4VnVGE
mKOO3DIZW6XtQiOczYL6dH9kKj3LxDrd/bjbCP89ClP93OmEGaaUwxQajfe4XhrsCgCdQFu51+Es
MV4a9tLivJv702wpMFlsW+XDL+odmbdew2PmGi4fMEnCbmoWkZ8/+64YgO9k9kuK+tTxeUmtARKq
CSBymgGGSDhp74FHJqN7JZJWyKrkkEWb8Rusn08EDyjnnFwUMYz91hpNau7cVTv/vCgxDdE1yTmb
It5cavKPuAJP2vbv4tXy96jy1N8f5IXdqrM6STDzv7M5iU05Hl53nw/pIvMP2OA7xCxqM6t4O4VD
0Zb60TDtG8rywUpLnWNIwRCvVFUV9BGji3iZ1+uJSauJ18suMDkHgOjBcIvFbWTTV6qy8LOoPA6F
MClosLdbbHR4VyY21kMO3J/GLeU1LciVZUwAl1tVUkak5xIDDH4Ucuz+sDt8ooQrI/6SM9W6cy2/
kwX9BhSt+WHrKxjQcYT1uvcfZmi/jF5YS82KfxKSwxDOULGMo2yrwLhFEdCPaDWGUmf084hdokZ2
2W04IynbqE2AIGCqsJxJP+9lSlBh/v8Mfhs6Nc3J4BNZBroBAbDtnSgIzYdVy/qcStPJ5H0RFWFP
KyknTgwSMavQyNSMay+j5SPgXrRXbVvC0rxTo4kEIXoWsiQCSH6wrRzVdhZ4mnBVDpS6JI/7ccPS
XllHJLg1APaDaeHhRs3sr5F7p12le6w7XuNdiYcCTMufSIt00PFeLbrjSMrf5eRstllYycdTugyU
sud/pFTGCCZIe821Q/fuWfgA+gNke7a3+PDzQdKWjQ/oc6guAium3a2lk/b7qO6LrGiIZuZhyB5o
3B3nF3/URumtuU1LWo82ZfI3qKn/jACzpt/MxP94bYSiW86twQ3wGx10CQl2OkPdcV8NPIslEegz
geTF7yigIZY28nmv0TdVR90NpezNdjokVv9iTtHHEvalylhrEiJV44p9X79kFxK6h8EGL2nsSu9f
GidQwEognvE7TDSabo18nFNGSSF5IpvSsmumsAFfHlpoizyKwLvNdatMGiqDUjDUsZbniSppuBs0
CVMjzv6QBCEy5gsUbxjp2ZYiq+gCLUyidXZyHQELrwiMWJy90O5WuYPAmHzskizPSWcztS2PbM1z
pt0GIx0N9vOonSlwedFT4ULPvIJqpBUWp+tQGt4IQjoxWll6CHHI7Iwq0c1afaswN2mgRa488iNe
71AFEj93jvVtOH30RDd8TCrYFh08wLG+sLDNoib8KFzoiWA8U05DvcidDI8dJiuj006bpYLzz2tK
WtRs412GDtGD/J7fCRSyvCk0qebGKmhjtR+yAqkztlb3FNzU2GtEM29+nJ1+AsxJxI4zqBo6O75g
EPez+TaWMr/+g0OWKQaW4OsKIVA/xN82vupny7E00Cw8tSbNzVjjif9svP/ABOn3TVEJTXpoxHU1
C7yj9dodPioBWTJdflw97COJsSaZaYl0qHzEM+5mXgEPmprEVFLsjiJ4IJby8cTKuLpFnXftNzmd
JfHNfzbjAT9rUvXe/pf8wW+s3ri1aN6RZ14pM6rPlrH4erobYoJ1Xhyo7cRYBZNpe09yHrVD+it0
Ny7Z/GY7S4cryiz38e/RTSwTH7uCZwU/OU6TAcpFWnm4Qb7vEoWo89kqbjgv7VlkOYuO/LbCB1rt
tPpuJwfMPkW/JpntvPaZZrRCbAauRUiCYWUvJHdOdODSbdv7nWXHvZaIRG95nZJDt/gdFkxYOaW4
6GAYnvMwtoDgyJuTcnfuegypjwAPoBR3oKF+sCmaTtkPTPqReveq52CP5dm4QnynWWCLKKdkv4/V
8QDSgEltd5wq6pvZ054r5ySJz3x0PMZNUfAb/UaxK0itaQrsp/IOq0M1gIZhVvWDHq479L1mGOYI
mbHczzuou7H4bVVjssSmgbBDkH5iZnt8uajDP5aDhcgZmLFz99+S7YMbV6MbygRug5Cz3DbveNb5
ounKT6bU8Ny+RoJJ9aA1d1fpi0LtHQtLokgely5BQlyzOntNTLlDQKR9awDSDF62uZ9XA6njwSBl
TQaqZlr4AA5y/JOxZgkoD0XM0VaGJTGSpkGsxIDYvSrDycX2R1FrR66y5rN+S4nPYUnAPHL08VC0
Qmpn0Gm7dhh+8nEPL8NUioxYRv3WRaWrc4BNkYQ4v1pK5zXsXgJ64VGtxpg3/t2LzvVs6Dv1aI21
z0Po3W3F1L9x5UasOivnKObymmaIljcGcDI7TAPZEuHpLVIcNSE2EL8L3gulDCuoK5D+c2X0IBtH
vGlZESMuvw9sfSxfmUU5wM5zuYGuK2x0esQcfeu2qH59vu2Sf9qX4es/+Q5FB5/1JBZkg66DN94u
Pl6PCgsL9FugYFzNTJX+B3eDqjGBHd47hCn/BEkxRSBLhtt6DmKU2/tLgJTX3ke9aFbLeCdKWY29
VyhrsFV3FkiltKxS28ysS+Av0xvxfqUXRjx8lL5Q8DUqMVjvZzztsaVv8ah8H1qC0svz+tuJ4aiR
uO4E4WRwII1T9soDF0hphmqseUdtW1W4RfdqljH3ZgiIYHGpX0DD6STvTrJ9j/7AozYsC9PIJzHw
FMCWCY9KGjfGG2ROV2qPjFpLIL5YohA6JV7kyIDomAoVuKag6vZthsaNhCXYCK51f0SmOA/PaoY7
7UZwzqPTNVoQQSGj8q/RtzED90b8lxdvLPBoS1fmS99ZCkSNnw7g7VPs/ROueIgpgeLN767BCjRw
E2St7tbFT3sF4iMZ3TC4r8t/3SPHp7GPxVvYEdtN2xP9JN4rKiMPFqZperKf2RRL5N3VCsJxBaLA
SnwbTpKeZSzmmdpQf+ZuWD3nJw6MBFTYzuwjqf3aznQW0VXh/1wcgtCE/p5FoiNAXmfZA3k/vNSy
eZRj8q45RcBAJogATsbaCl06OpnMjZhGb3PhMUnE5NHxErBSDQ2n51wpPATZZHMjdshtzml9WGXe
XnAuqf7Mz1+Qj3OKIo7uUvQN7LrGDZLEH7Yi+AmoNglvu6oj14Dqxya0qnKPTA8dcf7y7CcjMnhW
jnU+sdO6OSMkc80Mbnn4NHTnFNz/JA9yTKT4gLuo1hYQsy8ucKcckvQByJ0tAcQWme7DtdDhjk8Y
ZWnnTQpURk2gDy3qbTHGtPexz7yeajnxS5+MLbCVYPw7VDSsaJABz84poYRORPyVQ+ojw1Q/PdQR
wGAz+KYTaTQj8kTNrepIcEo4HuleDdRQuL1a6v2SExPrZQ1aiukpPeyh9Wt4jLBysB40dXfn2HkI
mZWCLYA3bBwcevAw6hD2x+k38PzfNZjRJkADpi6XEYVc5hWzSQFgEcENaTY4jWRSLFl6565+JMVh
++ENhJ+JsqSK+N5kP7lYq+4HOzdGrKJgJT7z/qlt7swC2ijQJ8w8Cq7ort0yohL66Yd+Um4isDD8
Z/ZZpqLa0jPxnl+Z1/HgVNjZd9HrJRCuV+6jcNYqVZ6c9UnVPu/eJj2Epd9j1GBtsRy7AFZou0kt
2GdPYrIag56Tf9oRWspo+ngWSMNWu37+dzjq9OWenF8fWjFdYxIYTPR2B2LLEPNPHk72KTz+lwD0
JPjdsM12aUAPR3tgckG6BYd95h5Kd7vrwDFP2QXjuSMWYs8A7kXBzKZjt5lj9c3SCHz2Lfa5Xep5
wj3RGC78c2FPYVCquFvf3y8+brzhoWiTayGOz4JVOh4nMMK9JkJPoveoIAtgkv/UwWW4fFfWko95
RJeRYghwJoxYAaZDcYdnjzmut2r+tNFnXjumkmC+ewUqqZLiS3xo9FRprnniMY3SUCEKmdXylKwr
SDXh/dSg6n34yJ3bWLnxhVwNMNl+ik0sFjErHy6jcH1tnqGkk99Ung+iTkf4krvgULdMHbTegg8N
7JQqCY3rWP/+W2g4nIYjvOrHin+661Fu2Z09FGYNdtO2z9gy+5Md1TbTkXfQWN0VQStWhVOWcVn0
jt1lPC5WwNHnWebkAgQ2rCnhq6uRWr9iNBCbfR0okuh2wDvSMmGGsq+EyVV8pxYxv1iGiwXR1Vba
nyPzTwu18pDa/EW/9jl+tFrxZiUOQI3dMEvezLEVDqZBhwPIYZdj8+EEADIUujD/zPtWzxhPdnqH
cG9brrWkoSx3bTF9VgLJr+03oFVbsvLInnAKwR6poYF+Vlpberb7KNHH9+r7mRl4uLGJEjPopoe4
7No/2RCxYzYpmr3Czyccohe7G4C5GKO3WFGCPDFW/sZc+/44lbPITUMlWpbMfMkCP/j2DHifqZPM
yAB9tetrA4A1Xc+WtuU9X09hTrhHKvvhvuyce+3u5Pc0CEiSMCtFGJvkNCmuuB5cbW094z1AmR9h
JOynSkiTMmuUJZ6iwcwXJmuGMsjReb0lj4npDMoJOavZItmrZTtuVGfvBhr6hb4vHzOYWJiTv5yS
qLbAjMX9Suf/BIVDpwDSd08p2UqBjltLbZyQq3l7ge5p35cUHYmEDKczrRTK9BsMrWSaCGZ80geG
txoPir4Tw5JijacMRbNZwkJnvwDOF6uGTfskHC+jjzbd4l76IH8Gd8vv8GYY/YFnmF3MpLkof/wu
OMgesxPPtEE+aOp/tXQ2ZErKMxGgWitDFixHeO8nUvDPqvZk7pM5QtBsm3pwXG5mO76+9FI4DnYR
e7UnyNdQojOSO34z216vAoPphfex8oRk/crQ/YYWDiVOVbP3GOlqehBAIGcXeAGC1ZxFEJXm+sEy
VrAIIkqTW/fAeS+2LldQzcP3QiAXspWMrIPZ7goLVzHJuxnfbuaXwWUMH4XHXsdbvG/pbvuR3gZu
MzvXjRjM06j8QK4PL0I/6QCImlhhxROBGBthtaz4gXD2eKRl9z9q4alh4Pe8phPbNzMD6n4W0M+6
cV4QVAsYrf5iogr+YjAwd/1nBPPzezRqo2EComqT6xxlXoJtg2DXqVMX3RMDEP19DbtvWNuG7NI7
nZ6THpLbNKCZZASN21YscuUKJBErHOzzflezSjxVKElivOwIgG2SKj+fXCP7/h0CUgOIbon524KB
3TgKXw/eOWOp124ynOXt5nMmOc4iAHGL7kKuj/pJAKVBTz41q8B6OflI2O5a/YJcTx2oXOj+aM4v
ovvsyY2SWRxk0dLk76tMFJ631m/a1gsgv52G+6wHkUFAzguY59hzkXcgVrx3N3vRAnWuIKt5m86C
fT0xnaEqe0v5rhu1x4ab+FoAEnGtS5SZyFAvbGAlKDO54skRaEXMV0GnLT+Npr/VA8vOLOERV1Xy
9bHE8sM/nYjk04ljFgjmOCHN5ZauILDLgWX+pVgCknVD7Dd1Yd7nYSx01M6ZKo0eM/TfQrViInUz
2rrDE9LdKgqOiBCY71knjYVMgrHmFsnLXhZnzXxX128dULMvnHXPYTCFoyj5UQ3b5PG+bJRrj8w/
W9Hj4gdLLoIUUrKLWuGR/H6tCzOzgcd/XwsSpyn+SD8mTTZekZGD6JsYRWY9SJTqLxqiiBc0rBlu
UhbWSgXbuEW7TzmEpd+fyndm/X6c3lB42ButE3wD2dzyYy8frDWSAlJdGWsyaZyar3xDk+cU2RhT
FD4+OS8AcKILm3ciS5/1RxIa6IbqcVtonYgywYIJLXkbU4lSU5McU4qJRgN9eP/SHUTpZiKXUUNP
ZBDffLB1JXzlB+GWHaYQjlFlazizP/d7zFLdrQOtjfp5efvLmLTtB05ih5eXU6JHFoljNCOmMawR
fhR+uzxtiYy88yQF8BHF+UU8NWhrawIjXcGIo80LT/n1MAoOrfP+KhaIxAm3xvEmArZdeAcOMYD/
4g7s2XmMxbYIng/oNrm2mxBMVq6Qb5UNatmqVDA2Cy54NTvgzIJYUrqom1X3JBgDOVWuJ/a11Ttd
d4pYePjgjpAv6q43/I4rUQUpruCfbZjmTIgbqj1f7UH8zpRTwxbgyVhPaW4gwelQVu6tnIrghCdQ
tavVIudev40eTM3BkvPGFWzvDcD68KriKghyjhhnWxR/AfblpYTBzEc7ZE0UNoT0pHGtZtoZDKz9
Q6cIhgd548D9LdWCp5oCDH5WHw8hYMTJaa39FYWoBn4g7LSvD7tLVgeO18pf9XPsJslWqjKR5ZoA
1CWnYeS76OEXDxNWT1DT30bLYsIEgor7rwWTbpqkPz4CUas4C465R7YkcglU3xAwhFF/hzBopsrC
cuUd4n54NXdfyTyU2N2EOjKegi/rFjo1TDxvll550CCruVoV/8aQqxZ2VbNANox6OrrWPsRHHkDt
hiAbZ7R2xxvN8UlGf1spGhoAJMakU7uTuJ6bqZiNaf+kkXvtGqOxwd0t8kh1CkxhbGDfwLATAUqQ
lNLaCBpPKF2rhzc49E4uSWxgnvyyhsiei9fI4tUbl4v9zYIBW5tRk1HeK6bOgfPn11Y8w8ED+1dH
XhHHUQQydGQIaVrmC7UOpTTBb20ODtmMqqL90pSqs0yXnzuLMVRZPd9jkbuqYZXEBGAFecu7TKSV
+LDQi/rYwhBSOrwOIWwByh8Wvm5Ygdsvt+fFGD4GNPGZWEaG8Q7Hy7LOF8Gq7r8R4diZh47BT9RV
SvlNv5mfHOD51wfOdcgWURbnFqLT/RBmxeR7m9si6p4wrywBz+Z/UEmD+Jr89AG6MaCwK5Qw+ylv
hgXvAwldTtEhWyweqnhWeup5evfQesEgqJK+cUqmerkKdsaFliuvaEwsOVRSVzPOdrzPcymWFCG0
maMymmSZSJYM9r3caeXCCGEmDFIfVX7G0jGVUN9UzYRBls1kNGbrCQR0ST+vox1W5srdgSf35FbY
n0Yk/9tw+bCBgLB0Gn404zJF3kxhdkC+0ogLmG5zCouJwa16KgKTeVVlL5X/vukLM32TViB7zuIh
moZNAzv0IdBWcAlrFRJYkyIccntonJwS7dWX1pw7Q2pnyDHurQ2zIa7kYXJgzQNQwb9vtE3LWypy
tPaEN7R5swX1Unz9WhM1bYR82ih/IEdGplqjY7qkzaRjdAEMwhvIPy1pneiteoZALpJeiUTvu86s
nk6GGaxiQDxE9y7mlSiHtmMdx8/MnIsV09MpwiPoR57wXqTx/C857yPAYevZBOpwP/Qdm0TKZc4I
2z9SPhK71ZqkdI7+LBjIQnVeYdFkGSnfYlJKjZ03HCcjEEQ1cmV8aBmRtZkBWak48FVhiwTI9805
IuW8PDU+d2egBmoKYkns62tvdpYQsAY23L90OJ12R6t++LeDYPc87MqM3CB11sfA/KtKvy/D2pWq
5eOBLzRx2Jq4Zm3Ol9+T/tWE3eLNrRc0SU768HmBxjYVgXzjZ9fK/YH2t/LageQ8MJ6JNozz7K0A
FwWlC/+tceyCWcLpin5yK0/jzC3jy9aKt6a/gVaHFd3qIUDnMqSMlcnM6rEJpim8DSk3TWK3ZDft
gAstTRn9bulwZmWAGFuUOgK753CXOkmW+AI+xfn0baucyxDW91PsyB42IekqGYBiRjDWCa7TsZ5r
xY7JInVncHjvzv+7zQaPH6AS3ZHbwbsrVAj4fEV+4+Vty2Huc2UJ+LJPAIglyYWXXYSTZ9u8u1jd
11EgwTddQBwvoPUo1Eu+CMjWXfJab/eeRchnIxsUOiE/L3IZ0yzzKd8LMf25DFMLUIrrzBaPZ2t4
U6tl2qeW+nCR39EJowcntpe3T/Bl7/GEhXy9hVM/xo92eT5DMLcp0MDekow/tW6PMgUzrMx06x8u
1LR/Dza5KOiGAp4z+UdKfxg8h/Ng/fWWi2f/EPwJ2jrNZLsDpTVEjM8Hu8EbYcVEg0buiyMF+xdG
nDsxxFlDtKX2Uc/pL6QPRsJwy4mh54KvcY2EAioS99iDgN15Dz/i26aWglhYUA6xTo4WcoDmaALN
aq7puL62U0jPIWBGHLrd2yJABNlO0aG6V9EkQxeEG8bHPA01+0jG3DcUYJnrn0EOg1wH2WP8oAcn
bo/zN0/HvPaO2o7GRb0DNn5naEsdJ0BRoZkGyCBXVV0ybl/rARGLPAeSjB4Hw8WVy6MAiFfgY+0P
Ctk2BT/2OTMtllsFHBZycR4OUYfbRmf6mfUw/KLKSJMlV+x5owGpXC03hjhLWGbhCIKAuammSmig
OecaV631wJ8/hNsMe3tP859UeCKkXSnk36gG04QNGX3bj+mLoLIAwT+1Ynb75F3CqO8/mP0RJk+I
P5wRSK8RAiX1PiLNrhVrMyfLR+XLqqwQLVT+4p4GBFdNI1rZE3revGvGDcpxHWfjY+KF4r/hK0LF
5bwuwNgV3yVQvFQintIV/F62H/8TGGK02Y0dfbmd3jRdXKeLpxMUsf2LHKtNZn1kBsfG1VbHC1Ld
02l82tdcnuBRIoEhRROS/nFpXh6UVb7p8jT5p2y9Rr4F6JxXX7lBdw/P7jW3tKFbJ4b6oMl0RgUu
+ca+mspptKnmvSDxMNIR3IJ4rvpIiyTagAFd1iYpfA/cDfwrDdrPMwt+LEofljqvtnxPSqEt4orp
WZm5iCRvAjSNRdBHWO/egra8dqAzScy2OQ46rz3GD5Nh6sa6PZx/iLxg4tZnflVQruev+BZGEvag
gKhU2EGblXSQtlZqn6V5f9Axvi6vkyaH5cKYAQ/Mj/0byHCUskhDSnrn7s2e2Tf8M+LKIBf6h2op
3doPH658exJGzXqsoO6vUvcQ7Xslcz+4kU1bqdqp8nR3/Uks6eNvbecJdo+qPsxv+3fnAufwsP4h
tIHnJA4iC/N7w7v1CC6vgQsnmSq7AR7HZ/to4SOfL/yHf5ukmb2XGWkUNHkJrfmHxFQtaseK2hHi
HnStNVDTy9OiWnUdiXZ/xmdbQMr7+yhpPUKB96fbAPeemovC6sOMSaKgqPHjcEnbbeiEdwz3nNhe
XgjmrioerGWYiDyxUwWDg3N8pbcLaYstlprsLUr9Z8B1GMiz2A+2jr163RBQPfG/vuOMH4M0l3ge
sD9uatCCMH04N8myvjtd03geFmOUzflgKYLBTeAxqHCGhuyzqNOzP2tPEdE4dw5fTgRRsG6mAKUN
obJ1bNxiDJb9WV0ptPgP82s7FZZ9B+jqI5qDHa88ohhtANWHjFLUwUxuYReQGK1ZCnWXgEB++0L4
sEt9oo9dx8AuiNzs4Rii8wqPM3/2G2TDHFqvWDDKXqhp8hPMkUvUH3lkXCdyn45TbgtWnAlFNIP1
Ybc9blbB8AhPI8+Kq+cxunxgLJDwM6bGNm1jfkWwTptqg7C+EvLZOb5wEer9uVlWyUjff/NKeItY
lGPFxGS63b6KpNAktdyDFV3nmu/grICamiXe9XsO8yphXHnZXLCYJrkHxBoIEF1MWLTpVMvD2ddn
aHL5QO+FCTK4/2Ly4/QL3a9T+HMtz0L44khbubgFIVj/KmvbWDjteZQFqLX6wM62+9NV+y55ZF/D
3ZT9RS8PXEmY1901IzwSsDkvlTSaj8wfgvZ70RwKiqPR8ZjzPWUcwBCV1XkICOL2q1mv4TG+kBMr
OS9dlFBQc9iX1uyTN2Y1ATFtLvMHBSW6/Sw0iiy+xH/YPHyPZ7VA5oViLABmyDjCmxE5iVXUDjjU
rLK7ZbS/srPw+OJ2dp9FI+6AxwiMvMnPNLI31nmqa/B2FJflK8i7nlJN4r0ZwzvF/j6a+y3UFL2c
pIIb68Nyu05aRkqWGJU5k2Df2EDcNaNzHVwuY451bxOjHtLRdi4LPRAN3sn1XgiLRc8I2SX+9Pc1
XGuyBdKnRSoHAYoPWijjcB8YDT9pQ9UcvUkY9bw3LQ7Bk6jvZdQQh5DgZK+rw5ggkyTX/BHBWq+J
71D4frooxOjNSqbYXe0QgaQvcyv4i/vxwVW9AxOsX+OfbTf1NdIm+S+kAeaPAJsT65Z+5/tnM5XK
iF26cY/8q7eDYnWvZ7o8dMoFc1/50Nxy+cwq/bkbEOFi6YHmsxKEbhf5Cpj/oZ/eRXn8ZtbUABg9
nqIPKqTaejwr2echMw5sSaCzbiComRKdFPNqDkgoHdQnaIrpg3REcFpozCWO7t6DEa/kCKmaSDrQ
/zkDgID4BsoaH75Q0Mlzgy4kq3ZDv/LFUgx5AiE+hGFaDX4Gh4C6/sF9ShfXrQMyJdgWtFTEhMaw
5rfdEEoLfGEDKw5y5VHFdLsovnGfL1jeBiDyqIzA7vF/EGZLypmL2Eo0I8AHtfX0T6f1BsL4wGFp
HPOWCqZZj6AynqD/0O3xj9Z7HFcK9Xh64vBcmkPYjbU55pgfrOoLDlYyRczZNZ8mdOJFrFmbZIxk
lH71Aq0js7Klzp6QnCdhODYTocF9UDdx/JONokcXXu1P0Euwbo9Wpo+Toki3848tWtyxjrD/pxxJ
2sfwHBZrRO7rCw8LjmKyo5nkGRdX3ypT4bEtdkMYp+90LybFud1ykn53T1w+EaXKQAI+YhWfTa3g
+t9Qhb7rfc/bsnIqYc5gSHosfE6XNXBzNCFeHNyMd7OpU0OyVScWPu0wM/im2Wq6/wLYUYnc6KMM
MyR0GKLVOO1oB1Nkpn9eTjG/BWFyFyv38a/zOI5XFpIb69s4MvpJ/z1/KT4rtiI/CgczU4LOcxh5
KjajfFQ4sdCM52OATsr4mLl7cBax3fQcg7Sp7BFvLSAnA5hpDuGDZ+/m4rGb5ac1arSC8Pyhs8wJ
ff1jdQnn8arFvVH4WsCoFzm0Lxa4tCXJVDU06T4S1z+HQIO/r8PZ2/nsutX6c2WM1RtDzj/kjqTD
7VndlgKrJOdHHKEb3MRNDg4hPm96cakfnb4aEY2VGo7wIpaG87RcqIpfNnKZnLY361EmEXcKriW9
tyEwX5jj8YHtKelcz9lpF2mOA7lV8b9WufETJYx6kC8A3lR25r00vTWBM2bp+KZxKSvZp4YH5d+V
bWbgzQZvfmsDbMUdlkQEYXN6eeZJFkwRdCIuJNJjghfxqH0J8Nsq58t4GoEP38uAO37Uj1wB8dS6
s6DFMREUgpO7rkBEf6Ef4Ur3F08mnr1Ir5ZuG9DJnn/gHce2eQ6cFy5/JO8lEEfaWCIWQfPp/WK8
Tvyfdk6gVJ14g8KaC1LV17qI4JCbNGjsDoR494FVyFodvajoIeG1K1unOzChfmhV26Q+gMywb6jt
+UWu0foKklsYWVuLjOD/2qikwFlgL8/C9P6GXOT7RZgjmiHFNkBcuZE0nGjz4S4iNYw3nGA0/uBv
hUbEtaGndrocbcNq3SCfK2iTfL3asOLCPqlWQH5Yz4WgZw6KZvFibDfgl76So8YJFHlNNUgj1sRn
DgIQz5dg7e489babecJNp/W5xffKxMeBtS09jdY+EDxFglwJwE8x/PbVDFoxevtGS9dhdjySM5zN
Mrph8Xm37UsJe1b0NWaSmfnyhieTmqx133c9ShDFrHiW7fr9h1CkRANfKdxaW6chfV2M5O1+HopJ
qswgW5HhxlzX32fGOCZfG8h/Qld+sE/pQxXonv3hyHc+Rw2426wd6ravba+MIjmT0dMR7ZXhc+8A
sov9+WYZv9VaweEXJFJIJNqikVRBtZ+nIvTGzH+g/t8M9OWJrVy0HJwcPo6399ckwfTc8a9IRBLC
q2jS350JQ0dGgbcS6Z9qojy60MUfaKNNJyDeACA3LcAvH/0geTIJyb8b7raCF6hJQZj+NXLoF98c
GDdWy8DynTAo/3qi/IySNxM9Wf2H/bQrpt+0Mj/Ys+dLvnhCkHnm/sgoQnyCo3JDnHuGQLusEC2p
aTKfEf5cz6OYbjwB+MMk15Wo7vnnyaq2AA3kyhqRNKZoyKoyOm5yY/ViROr5ehXeiuXkyhTpGf2D
RaeeHSf2zbl8F+yOTaqNq+aZJS4ElCTBeeQCMPv3oUSkcvrrHjBVugWWMaqFM7mtMVSglA9N6cQM
75HSrRkj11JpMQBF72YfqHOu90njdTjRnlqLUqHIodaIo2B6zqi+JhXyijZgeUOaujeknzwoSRlH
Q2byjNZLShN65jJokOrxXorbeKTvmGLfJpFKqDec7VNSKXc/1k/NyTvI3w2Lx5A7UZGWoZWUN8ov
8Idj/sb/fQtJcTWHtAcZhlyVMicCbFgsdZrMxnQ9owtLrHm7hX304zSaO6Ds2tE/7CZlXT/ShSYK
6w+PdzM5WHHg0LRbq4CbIMCDiemXjVQkS5N3elcsCYI3HCLL5CW72jsA1x5zv1JHDqpBLv9Kt1ZC
/Slx+Wv2n+KN4kQbVkoy2P5aNUD8v68Jc2u+7XwqhsxuVrj6wwEm4jiUxZAPBIMYI7y4T0smBOkE
h0oBdSqvteuDdg2LWjajrx8I5I+JcEBkTZ424kGrKiEVESLUbrodO0rGJTXTLY/ZFWHJJO142tUx
SefJiLTfKhFwZ7IwIMmZA5PF0bKM8FNMYFSBneqjdxpvkzA663HgIZC71m8GZ8TIYib1fY4niOpK
WDTQWGJxgukBQRo71DA++fwj5b4LdgPMdF5h9yvOaBiQWQ6OeIHB5+Tvtf/zCHao26iXFp6zjG7B
DHQlx5MXTt8DY8hstFjHoKPbiSlH24Yh16ubt3ovv86IkDQ8MJgMKF4wAkc5pYpA1Xrd8XF/23qm
Gwnus5hy0tJgYXMNE4Gz1luIbMoEExMlXnOGpkPK7+NRpbLS2tDzELniruMRqt0erkGsjwLdZ6As
j56N96pN6eifhqmHNH3P838QwBH9Sc0OFBlFVPciEnbfGo11/E31wl4XA1AP9SKhbQ40HgodqhXe
l7zUgHZy7wdRoW0fw3qQ1Su1zUTWWJZVpSaYDevpL6as9crM9ZisVTtbJAmMGhk3evYQ1xc9FcJw
G54CbX6Z8/4+yQChsd9qnEjmc+eKahocvgYLwK845E+AYe0Px4afnbgNMy7oDOmjGRhh4Nd6hBR7
FXSpV/Hj7Y7cpnXq/0p8MnFcpJrVZSLgRWi4871QWiRj/fUwJFbE8VLOcrOTLQzGFHqt4lCKiBJQ
AoCovRkqShrZBjejivhBj6qiJtyJIPikOTAiysPbIfcJ6xzfRriOzbD1dS/woFL3UNrGlt/Qwcrl
IM7+CotAMjE8YEZTxtW4cuUXItrmP4kgDRTEO/TL9iIknvSFmJTi55b4emW57rokVehUJMqgmpYF
6Vp8oRJVBCzImXsTVm8aFZV8bvSGeMvHkITPQnMyuGds0e1BZdAkgdwshpYqn/VmEL1Kmjb9BuZU
YxnQinAp3Afi5diyOzS5ejjDySKw8+VHnlTbqaO3rZgDXZgMg5lfzY0T510EzOnzLYo9O0PC3EWc
bELtYgWi5/92LQezDX2rfpzqf/p1PgFdM4teoOVddlb7GDFN7NAxqeq/Kkcib7AcBC7AOmYs5v+U
aIxfFV2e7+6ihxiYNz37rrXcLDOYw/QV2/x57YX1ZYAde6qhxoKL14g/IeL6AgJ0Q6wHN+mHW2k2
HEhXOznQ99gKYBfZTio1XAdE2XbNWUgots1p4+aWDe8WpPZvNNxMXDmqPCXeJKeJFfEdFygiDDcf
Xau/uSZZSql49XGO5JCnxNlqlCNduImH34nDZC2mdDWK3wq5TsXN1tCl/yNGoUTD3sOE0ARswqaC
ya/JSRboa3s+KpPZAm0BfkyVxhrLlDNMMNXQ3m//vo6jB13FAQtgY5Fs62/ChlTR9YRTj995iDqo
h/Kv72ZjwjRzGHPB0fJ8eW67E+n/2dYpuKR6Nvh9Skyi4eg+USQxbt0oCQMagIK5U5Tj9aAA9ZQx
OfZjpBN/mzTrIBiLeKzVMY6Ud/rI1N+KDUSsqk/WSlQxjav47rIehQa09HuWC8twMVi9GQtMeuNZ
xxco+HIPQrbOn1mx1N8bQwY0nDOY4AKnmPuvIebySiaNdkQ3FBQ/j/dW02akCtQ51NUuJYcnmUjA
O5NBgU2X9+wV28V4bSdE8f4wAgynSeaAHjLsHUgG+VxYsgmpvkRWUWbFurLLLFE24v4pblCNGiKK
HUTxIiiL7XXiHXhMnvXfv/oHAAUZqO4zqNDlb4UP7Wg8UrCOMo4MYpT9Fy8hIVNqf0nSJHH9CoQs
7yeYHA1l9QOx1WzuJgYABGjGLdXDMfBXgmaKmBwkqIEnBP9clfTicdCQ04SN0i2qc5K7J56m/108
4VeklI74AN+SPFZJxddqXqeNOK7eXIqVQX0mekiDD/AsLb93q6LDuEixGgjwl6Pb7ScZzgYUVlp+
VGYCYTpMsRXVXzIXWObXqQ3U33c3nPt+gHsZELAL0+jTuio+rtuYXeJksqv5kxp22gnFqnhv0JDt
2nvZHHWn/gzPrITqazx7UuMGZQB9dJRTqx736exaKGWwSaW+BQVIWeB9t8k95nEkOZjlMBInFwPr
7uXwtvsO18d1MYHV206bDrfZsEeE7rT/M103bOdM/poFnVDZnxMzhvQwY8XW6A3B63VA10Q9goF1
rzzyF8Nh7wrAyWrYolTeeJef8EKXWDoREpMtGm1fJJPdjNlsxSl3fihcXz5fN9Hzrg10dbdhgfiB
Jc+RZAJh1MbdZi8DKiHQ/7MTdVCRg5jKh0/ifz6BpZNWKKh7RjCK4AhhDx+aQwU4tcVXXgJ9s9vC
NA41dZyOsY77wc8eAvVJB2Iw/RmxoUplI2qyZV4QqLjFJjV1Lk3FqupnaHDgVh0R6aDNxBKWVQ+3
s4cdEOM/WRLFNvUJbUYLIoxdK0N3dGHWLOqDb+x50VmHUhN7zBrvKLNp47Gq89LRVTXEYWCSl6Ud
t53HrJ5w4PBGgGY4RAdqIPHk5qjH1GsTM0Gel2vzbUuig7HmC9i/JxvIHJVsBy6VmcGGNAs2ihfV
GDTVXY1S20xI8w28zENSip+RYCTeiGuw0fg+AC843UNnAlxVrEYMxgSrU9kv8FLtYOPH8pXiZQhu
+fVF8BVZUqLV6sq3jEf0ZEIJAtZinjpPRDmPBexaoJVFvTQM3WXygcQpsy1r50pIacYgcU2VfFrs
T9SNEdtyW5Cesn0RkVZp1OG2qOdFGVPU2YQGW+0d3m2qkoxTRas4cChHpuIOALFgA98rI8viJKGk
N9UgDevAuqbKj2skc62xttBk7D8Jw5qtQ+y2+vsvxs5f/xjW/WTDBMZ8NW/UyEhnBDlZISFDSVYH
rQpX8uacnTHh2MA81IuUmkm+Y5Uu6FF2tI6YRmcCO5QfMJNyyxObUs8sPlqXcEKFYQznPqEkTrLE
/jpIlYx+l1e0qZn0O77b0VR7Wburn0h6vKLKGZD115DosmW/NuygslyU1G83UQ6zS6yh/GXxWGAJ
w4ZjWb0KhWL0EKYeGcDg92yRj56oHF4/+nqUwfyRO92donCmnFeqdGmgSi+WFbEtS9RwdtlYWD4u
uaSRSofxwcSkb1r1dh9MPI+kTrdMCLM27YE+kZgOTObIrMsvQJjI7KNvYOqqRnswSq5MSk/6tKcC
bj+PJuj8B7W0ib2O3R431x1BvuZ7D617wW3TxqglJTQxQdcI9L/41EJ9NjBINReEByPeBgSieoDH
OjhAmFnjnz9++jSRcCgXbhcObst8mUEVRtB6ibx4Vnf+w+9MKJJJH46QatcUcl1a+GktJRvGjCZS
KjqsiXiQawjc4i6YiUbscfbjfG1P9Fc1/hVhtbfyCHEtb7sKL4aLbVE8V8K8wMXpEYZ/4R1iLxPS
NLepzd09AhwVtEBcXGRs6eIS+9XvsuaVbTjAKIUJ1aHxsKjEwz33WWGI5hQv4ZYKqIA29BePi0c2
YWHWKuTzJh9vIH0RC7V5zNQyy0lPPkjfYNuFd0fnvmPee76NZ01nSHIpV7NbmCcY54OogE5vZvgQ
B4AiNBDpMHedHEfCQ/UhUGpV7kF43+PODVgOcMvcARB+Xh8DqXNJZuTXIut0f4gTrU+N/+1F8AL7
ETcQJVre5Sji2EusP8kUSJmCCbj37kZSj+0GMfh3gToaPYfTXzj/wq7ZIzmgXfYjipYHTYFLV4WE
5IKys7jx/FkpKS4N97ArjEFxDr1ZCzmINokDesmw3SGiGu1ZrSvE5Gh5fFIjPJc1s8pr9k5xCpi9
CMzNKB5iH4S9hStHTRQ8cyBlycLFQUuWGdLfQdzMlt70SJmqdCCKjmqv679bpEou7QGq6H2wmwzI
n5V7PVyrmljrzqm0eUuDiGE5c0So4me1y/uB/zfGCAFagkoH2ZrNI9vQcOReljXBnPsksFdXC4Dr
u8VVT5977ZE9P2S29junyvj7yuifu6bPNKGqybu73dnMh4Cl3NBWcP9QU16b0O9UuTyrOwyvqR/x
GlilKOlST/xXi2Njya/mXi6nPomjRCKn5seV0qy8O/Dn9+tl/5BBT64R5i2QVf1OKemdCv08sX/W
BqYrmZb/otZebwSLgr2QA0XNnDGnW/JPJvmfP6pdFtpYNEZGh+wzPAyc57YWDwF7MG73gV9NEu8p
KxPMPJ03z/plSoBwiXcCgdMlaavbUlAY9Ec811CXxXbaA0QtJ9FAY4/w1TgH3bk2IxZDB0Jm3f70
YgAIdUfnC7+Y06R+x5jafOD40VU/ozKBZHkYbC0sqza9dmsWMprEud4z9EuYHirtbjxNYoXGZYUi
AEsI3jKu7D9GE2MMGk32p4VMgwKyRX9oXGtcIekKB8lNPvgvi6LtOY85mpJ3I+PMILea/0tE3uku
OdFx8wtUmB6LOzS7faIS6g4QFVsx6waw1dmDCx0kYlPrM4W41a+OeM49XCUOAcO4+H0utbN0dHM7
h9TISl0owK5IQHCO19XzYHJTL0a+INrZ5BjGf2vB5iKnlNAT3RPY5sOTRkoYtx2vrJHH1fwEdUhS
8XrUnYKaxF4Rl9iN1tjYP1JMuTYEwvTocJ/DnyJ95gYaDbhZMibWjRhgN1c2LbeFJtDoTFebyKSD
tqw3aEQLTFpSdFYLdEbgxHnlIjF3+nuNYrja2d9JzGc3PB0cgWK4+N2yllzwc6+e8Gx4WcJbLMqq
GNheROACs5UUApB8aZMMvMJa6EZGwstQFHoeimTGXDZmRO1LgcGtEBmZrMSWplh+0ctQyYJQcuuX
2ZaPNXpZdxGyp02gRJhyqJ3upmVQFSWVHUmRczlh154Egwc2UXCt2Y3hWcm5Hcf0O0c+8k2QB5hB
pWPaIVmtjqTyXAiaEUpxiZhAl+a42ubbCVo23A4dJeW+omY7qUtN7zkWm69yPhUwNPUrMXXWGqW4
59gH4xs5HGerw820mOKzh5L1Ux54n5disvO7f10VF1Jj9LswMyJ9nbtxHteyLVmXtX17KmcJql+7
FM5tWVgT+HSlfY69exQZRChiH6Kg9sVtafze1pWWhN4rKV1t0E73f4P2FI/LpmBkaiv3tcJe9RbV
t/JNpSapieudvqlIGE1CuPYowfqQV6ohY0zEoyoUq1WT6gP1onSaFTXrcaJxXbef2y3Ysd/OOZnM
p395ePBWzUD0OuYFcHJfbZa3vp6gR6r9fxpf+f23RIkYjcVBN/MqkfXP+pCqoryI7XjA/DKA5bnp
wcBGbJ9feopxbya74TcqwFarw9dBPfnfe7hChWR57MI5paYxJFZILsPEpOunlWBmyFz60KkIuol6
r8RFkL77J9T4jERKk4bGD9p29qA170bcfnl7pFpJUE7dBqwJmmm0FXbzCc3SawBErQIPq4aL4kQZ
6J9lvnk+iN7IK1QlziG4XAbIT3y42ANyzjT2nEHUa5ezJf5xxHT7lbprNjMMBcgtI73AYAH/PAKg
6d/6YeiK0dqRRwheSCWkAyyCK3M5FhH+XfpaIaxmUWWHYuS/c1a4oCeBpAtCIgwp0kgZHKtOlFLA
6wfYLFv6x/wF1WPszYx2VDsFNfR6RFdQvQjNgUBma53awFA1ER8l0Z1l8C/KamjmtiZmkVBjQQlV
3DJvsP+iKq3+wwm8mNQruu84i7GjaS+bvolBpiLeYiHonwM38ZFST5MB2drbbS7PV3k2yc0JyNgc
1AwmOO+rxHYb7SaUTflGO3imylqQIGxZzSP7HwR3i4uXu2TTe2Gfr0G+Vt3TEpZwmjbTpxPgTFaI
Jxcr3SQFv+9P1dYnZOOcLVdjhKmwE4M76HzexwvMUbYygpOVeW095MzG5ZZ4PgJmtme+AWkMd6wk
Tbit/xeFn/SD9CklGe++wDmKyJjs2hpYMq3Uq3cNB9Z9xB8Q13s0y9Q4n/keXa6rwCfKPNQIK5Ko
KfveLqTl0/glBU61sddaTxP/64JbGlQYKTE2gGarlC8G3tNcuIfxFSsorOuch9iwF9+t8JKt5lnH
Fjn5LnQEgD9wxURSAKykLG9/oHuywHzfJA8iEtLPxjNbv5lfWIM+dJruC2f104rC8/HXzyvX7G/6
zvPsX30q7UT3YWTw2hmWVHuHZfTyoj5Shn2hSaS/TfWWKiHh1JmmfdNVSe92YPwJfxGW0j/EPyYw
6crdlkp0/WOXa6KS0tF+NPbe+z8ZWrdcXjt2K92OnUAk/cshigiBdbyficxEB52pjwSenN7Sdcky
gxIizrtAPra6meIle4xuKpB19bopLs8IkOrSW6vojIjsCw+C2IpjdP2/BWJNirI9NAPlYI/czvYK
p88k9PjHIn9+2BAYtdkraNA+pws6y8C7Xzx+cqsioRCEMGwyduoqs7Jhr4+LTYfJ6FJIUg6MuoGg
ewKAfwgT1sHkxoMfprzmhoRm5G84IOrzbxc+M/CYb+6/IqdGbAk+TP1JyPfZ7GnojAYmnSeJpRK6
4QrrfcJlz9mT8B1NAilYmAMRlr9g4h0beA39W4MsPrVO8x82lHT/4Jo4k/EFHwVqr3GGevYT/4SU
10dMCTSxeJrLDEtZqwaFp3SNMjD+R07P6BTGQ/z+rg2ykmXxVeaCKVy5BI0xoSpgS9+cHh/khiPa
q4J0t6ZT4T311GGXN/tcrxf6UMcx8cL5pTL0AFxcN5wTgFUrzyL3vHe2enU69muyPbTJCOAvpiIE
y2etZs2v+yn9nYcUqqQ3nfiHr/UX0qi016IjD8MsxNepx7hX624NM88KcIofz5/dip155FI8xpFx
TQv2MIfFVNFOoinotCHAFkZ60J7MQ3FqXAa3l/Qy2RemlJok4ty0j6V58bJIT0dW8ByFF1ezodWt
LQJYo224XwlLnO9ZQNfjEgThKdCobnL8mZb999Uy2wOYyL9ZW0APS+yVoxuNgOfPqGoP7rOfQXCS
NQH63dtkTcRt/eIISW3g+TRF/6aISm6ET9weRpQkH+aVdv8Ac912rjJGEzq9cUEbztb7ptPr/Dye
DLQoO3ZmTbH2D0lE6fgsjRiL6S/Ly/vLbLyYqMS3FjN21nZNBptLzQRa9pS3ykdRghvalbFCKJ+S
gc0TubNpAFzWGqW7rkLM1QhDJrBy5MyRdl/PyVRNLTtXUDZ6fJftLRxVxj5LwmDXmJE/c2bVWYUI
TFNJo7SjmA3MjOalRd/kKtXlpqlwOWujsDIlOaEAKy+BucUVUXtWWc9qUK1vlrk8OMfZCgN9Ed+Z
CK0/F9x3PUOlF8gxYth6xDAuvIwvNR94U2GxRVvltcyT1TTGOC9NXKzoBuM3u4xzkEwgBAzha87W
SEqW9yO7xX124K/mzrAUFPN+1sXzv7k+nykd290UkBinpM+Pr4EBLgVASBAmbMAoGjzcEtB+Fwe9
oAb/NTDk9teto0khAatjoybazak9Qei3ZurM9YqdnTm8mlan6d2b7WfR5A5h5Jd3Ek1g1QrBTBFh
ZD5cSpQ0uLTvUWnDDYm+ITFEW9pjLENKa2NAD5GkpeHFmqsNUGC5xXHxbV/0fLtepZt8WinZ9JBY
/rKbAThDVSjDlVFwmLYfmqcj97fkxKosEsVq293tJuemd2wMoErCtg/DGXOaD2b+PgZ0lOUvpRgu
lSxU6ZM8VFdfY0MctcKWNMNVAij2keNd4nCz36EnD16t6pI2MJXp0eGrx79rnyiSk8ssCyOfPMnO
pPpf/fvc9fYcjcp7Xpw0ql56J7zWEmbjEgSrTYgl0Y18HyooBWJM/nMTW4RiyEU7KN7YKa/5SEB8
ZiqCZ4kb3dBO2bs4PZ3T8yxIeXJe+XlxGzVIHJExi3zekYfbQFgqGw8kQfys3fvbwN92G/CH59xu
HY6/3rZIkuDF/IvAwg2bdh7DAPCV3NECOXkYyGLr1aIT0bENM08U2efjL3ImMW0j4mHV6onnt7dr
jPev/d2AVjdFm+uUZUcjNAni5NMbcknqtKg8exRKTAdRGw2pZI/j/nt9W6+gbM18YniO2CtkzGPp
LrAtytCHqRRtAu573+yO8aK8EwXqCD7uj8qOv62Oo1wXTwBm2nzeo4JYpooJkaERnqMSEiP51c7n
iEjUC+C80WG8UiH+xapVgXIyLIMw78gLifvwWebmSCrEaYjKrBQvpsNzP5ygzx0Tlz2eSm2frv5u
EL43wus99YwGt6jFYhyGoe0Nu8uQQHn2++EVPVVtGgkjwrKk5FeE0ZqXSctFfSkAXjrbY67Kt6GP
8A4mlcMvFkScOc1Wr18fUcFmLbB6n00TgtaD4Ldgmn5YKqb9qPoh9OM2TKfcoknTu060vZQsEkYn
GQ6m/iT/ftp0gRZpVuRgpDOq19X+/3fPJVfBWIWjPjKMpHccp+18xr2rHHkAarMgJ/COGYpL0e0s
KEUTB3nFbNSto+TautnjbpQgpoO/LohJz/+MUQOHzNJKoz3/s9N6D7R2GoXjbgj7m2V49CYLeLHa
H893IV8Vk3x71BLY7rCtzu5MPZfKMhhQlG2oPxZ/+aShyT4MGWYCdhhHJl6UuLCCxBBrnxjVLbHg
aD7Pv/f+geRvxRR2ovPFBDbxKYMKVVTaENGRYnR9nkSFUdyq6YQQuBHJHrFbtJxQ6CAoj+Km/tFa
GIboDXyaHg/rWPWn+Dvl4ZhW4gCx03x8mWMsthfnoCKNE8prfsCF4VEfX1KcV0stniWOTMsvxxyG
5V53BR4VbaJ3/xAAnP6vBGMf/9K3Y83556TrjqNxg2lvMTqY0PVkg8Zk3/GTtBgNkV9XStUGbtJB
OtVL2cGgq1QUX/w+KcXibffJmysx7QTP5HGEZ65eRAhNWL8mw7Hd4tbaoTcUCIEnKSao3Z/ouXUO
AImxR+cOeqG8C0dviDE/l4neaAcTyAG/4kyZo7K4T2aP0/7aOvquytcGb78oUZv0nPZd4zIjLk0y
O+pUa31FZAKxvlFvMMna7xD1VsZhvbh9c4wllMkOgx+b8Pi7AbuWnqWR58nN0uHWQY2xnmKbsbpF
5d6yRWj7uf7EIu6/nOAMTCkAdcQf25JIn0PhVNZImyl6jL1HAmpLdDDFRqh9WQzMfROXmU9bBPp0
uRudDPtPEI98NhZHn2poP178Iaq9L6D5YOK+8Ja/IstBFbQVEuC1R5JW164YTnqtThj1/xfenBnl
rcQKMAAMadW0IS+UwjNpMYixApVOgpUcwejBqZitzo5I7ueSbVAO11Toh02JoykjdfN+hbqz0Z8O
HPFpMwMW8lvo9Lk1z5mdiy/QQwbJWB98n0M3sbsHA4MCzzcT9r79JmiLslWP+6Gn5zZbyzp37TaY
YSfM7jtO54DCSOVT+Ecc3D9EFVDPPjCpEK/xqpp70TvntLihDOz5x9QcdsdCDHBRR1dkoVWEz0Oy
+sjgF4OKqw5NqCDEUKR9pKl8RUbz9zfeXLbhQUOFZowpi001C2sX+K2Fpln0GJ4+tVuRpkDCrvGA
SvC77ooQZwJLVduNz0CWft3JioBpg1Mncpbs5Haq/kZ5qP89lNqyVHt/ef+EbSy4VOvxbGxS5d4H
kufp9OqwGQzuFbIN2qYxUPiZnVSB1JniCt3F5xBJU1CSeDxFPbVc0b4h7imu8FvSHs//FoHM7a/8
B1YFst+JLqaJbE2kS0vDIn36zhML8B0YENj5APBfEqJU02f9feamEi9BoT4UOca19E1tBuaXQCdX
QqwkQ8+CzXDPvQSMj7htR4qwbijAKVhoMM0bN5T7uPz1MObN4OATF0PmOzbrUK92wnTfYXPMVGhg
xjHv5Ycq/IkKL+XDI1c7dRMbuoGTB3rKc92kUo86njAsomiVGdOkh1KhMx4Vi5QPiVoE/pQXy38h
z3Sw2HosbQblI9HdxrQ6weQQiKI3ZjEXM1dit7rt76UMTIHlhquXYf05iJPOgqgVvEOKqnLSZmgI
hFPFNFDCpvsBX6idvYaVBLA/LSVp/OIzFfayeLf0GK8PnLhTZZe84kW6CtFQi/zA+GTcAaR9GHv8
5RfOPTKON+QN8wRc6SGMF9NTPxqb6XiT1AmwqTGLO/oLYW01eGz6sPbLJH8i1JAMGxFhmx2/agzY
d5eOAV2s0SBRyfgtzFEhWWVsM94qOpiVVuLaYS+cMk6yR8nlYnaIfRxVlpiMfffiw9HO+wOSJYCH
3OTITF0uj0Fh8P3UcuzxDkS+dOXhWQGf2G+38oWhKfL5MQMbj2k+tHTyzyANx5PoUQL6oQRwFhI+
Tsn+DcMpR68iKxS8PeMJOaEzlUady+x30Bq8o63nmL0UHdbM1G8Pw6t74bnAzSOLsVIb0zWGY7e3
51JnJsqEUUMhyyGmItV9dR5UvFMHwftIeY7rZmYmwsFyyJGQbeA6CRie96ifelSxQjFvCGGo9N2i
zgSBHdhixtKDSePnL8gB/N5s7hZYKcAd5pu6LwwcYUmlb6RcZ29vqJ6vv/EFxif8aK6rN/ikrahB
ZT0EjyMhLACc+nuf/vH1JRdCf7/7IJqOcU7vuEjhKuueW7E8OGQL/NCqGsNIsbVgHdNGr/Vs3lMc
2UO2tZgq7dnlIgLb4apOHNVX4SkNGLRLJez24OC1bG1wRcpdD+DVlioTkgdve1P/HZ6feHvxKJk2
O5Cj0KJ/iD0an93gpbyZa9lSUrCydfdOH/ZCOdEOS1pbwBmwmDpHSZlByVFJhpjh3ubvnS3VKCg4
LBENVhUVf5wY0aAXGbG6WqEqRBR47simjYgoa3FjMneLrrWAwAsuJsh0boohpg2Iec4e7MvmhaCf
hUhSz1vmTgfABh41YkMvgzvEb7uPvBoDpeOhC+rKAtjKexy+bQcMpgfXXILR3utqS0easmCIvQWF
+NVgJJnHmytj+01yvEh61Cd/6heKKtK2fX7WZVKPJtlYexw03L1vYWKD2oZOC4yDjm1yhadOwIP7
4RdeeG1ylkplEAmTXVVXF8JhEKXenxTiGOAyuoIkA9BqHu4XMLLuZCXq5YUMoMaCnbT1Cp4ihOqe
HMml7SjQErkJ0gPw2GKQZGPbi/goCB+Kr4ulcg0F1ByH1/13uzm649Lk+qQwRLplZhIa/hzkRaLv
LIw2RoCJcz/rU6erLI7Y7Tp7lZGxozOHqvhfd/mkF4LnliGedoljMbMcd7o1BFeHpq87IFoiI95i
L0m4M7QIQ1oG2d7fznq/MR0Qi5BajBzjjusywyDU2LuqASQZHkTKAphZVkRJv0sAuT1O0LkwXmte
nG7rwJ0v3+MKHOnnJqU4ooRWirMlbIVZgpQTmYjXNlFPGvn/utCZByomy1fRZtP3db8k9KhGSwps
0NvaQPJtZ7J4/yP6rtJ7/iZpO6ZARPPpQoL6th2x/I29SoPe0zCSS7X2e7KjFxzbIia1uMtCsKOY
9V5b/C11Kw1iT3fL13XAZ4Go23rcGY+ZBR7AMmWpiC8mJuKLw3O32IWzTvn6DJhO3b5ohKjA+0Oz
TrzFHujbP2uOKuoJUjGAF65ADeQ95gYnrvA7Ml7vQrRwWF0HlLdGcbX4aVvTKke+t+E47poOfr3M
qYT4BclNBYtb7NRw8ZRvC4WgCIxBfzLzan7Yj8Jm8FKDiIBZwwrJtecxSmOotClZC2yJ5xP412Ue
pQDeeEYrd6uPkrBAbsveAjpWZExtmiEDyl+pAPqnFeNtxpxhldNpJ3Lk5lEd8xixmgAlP8S/gl/b
4rKmQMlzvnhtvjt0CoxAHocVExUvWFLjuvW8k3mCN1iA7PzyMX1VV1dvvai47kqVsMACWxfvIc2F
cGHB6BCTqb48h6celkA55fGXJbNMjyGqK3GGS3g7a4vJX/a4oQXVr6xf3TVJ2pC19ld8c4ZDiwL+
Me2bzjQhH2y8vVpDuLIShubZKobBdRzjBj23pH3SOG7mmxXNJt/C+eM2AdmOV6F+xuWtCcKIaLa5
aN8bXI/PD5YfIIa4nLpaiLVRitAt0E3j6A6G375MH/m9MoIk8sxrh0J+U6+9Y7zELZMElk/wPdsc
0M+Cy5GAK9HoG5W9KiHQ1vkMy4u3S3D4AsuNnvNMfxWpdqone1yxQY15V5JuvRnpcKSzWNrn9IZT
CUp+1UwsAt0+YrDYyhytPzdGrww52DvmcW/3eKdZG8/eP6QPwOt1pjjlDQ+/ftKEjofkkN4SBrqq
Szx3hikbKaa7DwvhQQJeXIg57DGIeWdu0l/Y7E8QluPbdQDtB4K3MImYbDcl8dlKh43rDJFL/oVj
7uJALzQvcwL9v+MDwotOxdEsgcllzm2pgj9w4PGYv3857fDQ2oJ9FjgOCfUqYoSaqPZ58cvLQ02r
mF7sBdLL1pl1cEP0xvE4MfbRk7jyuhsfSx25Pf1kHmFOSiGk53bx9i91eQkr/rkfvVws0yd7WRy/
C7vRPgz+a9p/HN2czTH7RjePmCEgXHFIsvUcciSM5bsKc7Dr21wq7HPcA5QZlhd4ZLFWVUnoZehn
OedOQh+7FVThIWQIh6UNGewWoLCJ7i/VL85mcUheR/9VgqJzqMIRA7z5aZUaoTDVB6ZK3Ipolq1C
9BNjwhP/tVAxHxFUTuG0aY9i2+J/H2prxZpf9HU5otdXT8rqZn1H+oK3qGmkOk5DHrqDP97AP3pn
RFGkUPCdcy5PClrcQxKyTe3eFY2vnisc75XXgCAUA/qeQprJ+qMg792WpbBwCw+RMEZXbETCjlZ4
NVyCSOs66bRNOsTuCRkBK5ObSBub9/3p0kTP/sg6OAV22WsBAgcigyc0Gw7JauFU5d92qamD0NxZ
BO34KNRTRXV8dXBKJCOrGdLNjTPoLqD35wZUt1U+GAC3Kl8i6jRFVl0Zk68yg0vQuMasI7uJInKx
ykWnjRPvgsTt5M+4H7BbAnQazfaIT4eCdg5+5p/D35MnNcB+vOEu3uIfhP+m9IWPnnYoA5whftvg
E0DmuSY6hbo8cGQxff/mAjD0vQmkhPKndE3AfAREIsAJkGCoKnPTr7r5KfZ35sFHPLmfWK3908/0
a6sWmWay0Wq4dbrA+CI60F1UbG6TwPmAQEtnMnN5tHDrunvv1EkTbE6dDVK5RK5wqrh3x5u+g9IF
lvwI3OF2IrqutyR7nLSbMYccU0ZHupHfmEAJxith2zBPGoni/0ZbsZCyGA/uwSRbeWx5QFgcqOPy
6uPRkk1rsMjOMUi3MtY7KEkDToK9LqurweDvf1whghK9Saf70fb12v2IO/DKySwc2CTacuq8quk+
Bw4RYscBYfYS2i8uieTHan7G7GbLR3j63MganSKFpxzJIGR8H5evZbVejVZI4+ncirPQEVfUjsBA
LXr393qhrBrCAOypfb9i+T7n6jZBY6sYyMhh3rnj4jEbhvwlrQduCCR0aS/valZ57nYTERj3KFDi
KwEn3Y8TXKg7RJcqFIhYyqLPM7Nw1IhToW3hy35CvK4bU45oZYr9sdOCOhsrlWi34WE0970g/6e0
NZLxhy0oU3sDdOcOPwUI3SbwwAVDUSJEnKVw2Fs18kHDq7tX3Hs68ZQJXr5XPAn4vMUW3IBEEKnb
6dX0c3CC+X8rbM90YWVyucvbVKfY7saTCv+AGDxnrVn7Kr+45/pMwB08zEzPSicXue7Y850AaOjK
ewT9UMQ9ukE4mId+lVAYsAYmcljbuTg1WhcK3E/qxxnRfZhxuLE/5BUw5opjDKDLAqLNaHUASloT
Qgo49NN5bMLAyoTGyo2romPiIrpr2WmjkZxREijbTb45Ixwafd3cmDVgyR2U2aLOTYxh1Rhr6Bxn
/iqmr8jFVDqpRTaxpmG8AjFAPIvn49Ai09LA3vlupcBqKkk6rsu12KycyK9KakV/YsPT1uNKrF8d
45fEsJbce1brXX+JTeP4tE4VVO5nTOe/EVQHt84u0B25Y+COjkVkRvmH9jYZANxkyFHTLYfdE4lr
bievjdKnt6ffLjXAZ3PTEVCcfDRve+EsTO0r/PT6sYzPpf/gjG6jL4X3srpdP5s+MQzlfKciIQxb
LIuvLUN98hrP3KistjLvE6Vci52EJrOdhMPLKQwE50hjh0BrtoPojP3wCGulmU0WZKDwW9iafIFj
+FgxnYeH2HXNMAuLJ0fCV5IMyKLVnWxAYhetyQzei2OcjI2/Y4ebhItRp7xwTmtN+8U9anscguvc
39PMMMNzUH8z4YT7ILhvwlKtJBU04q0CacsO40U9//wQnvtKwrLKuAja/swo8yQ7losFt4+G9xXg
dfkX+uxZTTUZL+C7yciAA9RhMkLsY3rx1R8B3W5NHJU1cubsPxtQp+xVCPldniRDIaw5Aoixm5/g
aZLlfXzAmlYi+oCddMNUTp9ADTRUT1G1ejNKxga/kwQdyq1WE7pCjUj37cNbEDLUEDf22pFHMPNs
WbVTXG2EYkgeEOCvwzp3zNJ9j9V+1SL3/K2jCpSNNsyVLkXMgVNF2MWYrpARpIrN9VZsoc5lMV2C
XvcM/Xzz7cu40Tkri3Q2aKynodRHowX3q7BnqjX1LGfr4owFFELdj0oURJmV6bV405zvcjaj6tkh
V0Y476e1tWDd9xmcruvk4ZtgG7nTBdl6OEwS/F6enHpbRA0wU1CgDmKkxW7fU1mqGJ09Qc1q65Wr
/F3/1ps64/j5BTxWj7lfxF1EZiYFdihd7FLz64eTzjQQEk26BWbUHur+9M/lEVIorLRfoGwzQoyl
Udqo1p86Z2w40e7nGgZOf9k0atVvOYMNfL231WIa0pouHJydld7fWivC2EzA45JPmmDRvdrvqywZ
/EUPf4CFTbyHndpvImds/3Mh+hh4yE2eu6EORPfSwaHqtHyBtWyKBnQpyaGp8NLCEqPZaA5kiGu1
NgXfcn93IlAS9ATipFqmMUM9KoTpl+LH8/4BBKvtAzrTk5In2/pelQTRSmibh7pewUtBimek/kjc
zV4m19wGi8Cig2Xi4wHdbe75gohjW7hM+YPdzYoK0qVosDgi0lLMQ0tXKgHjM+MTkgUaJn4I7oTf
0oDRJcV+o5cdaKl4b2e1C253hgCioRxshp52RLWsKVusn2ssZjG1mn6daPKnvneVezsu1PYbd6dV
zauJSugNbbw5VymnyRXhpeU85DzAzaR7AXABbxLjloBjZNQIfvnNtXsQm4ToDveVC/j6+PwNNmJ7
hS3aKy4Erajn4CAxZG73jY1ByFvzEydV4BVadwPisiP32e2Ba0sOKCIHhorJSlzOft4JDeBfw2iD
y+/cb8PKGSblWhggeDGCxKoJYpdict6Z7El27O2/x/u1rWvlxy7jqc1e8MO6hFiNqB33Lm3sHrER
iGu6sfeFRhosk8no6WL0jS3U/YtS/O3d6gCkmxr+YO+LLWmL9wmcR671nISRPqbL95IZ5KBjITAT
Sz0tyUIgi02ccbM0jSv51Jo8j2Jo90Va51hSaK39LuRDyJyxsWdHG7f2KGKlo+qt1dAiwBxrA2VB
Gel4V86kAVGUY/BvuWsrrYLXqoMxaBBq/fEMX4su7lrGSlLBxXZoPlYgTWvSzyITC4Ny14BJ+9Ak
WhTpYMYgx06cUUQAR/SyJnxSSUSHEbuwyf99kJ5DFCkJQi2yRbLHlNhXqbzl4R4QP14g1da0/dMr
TbKAgOhDdqiA6om+tbyQLIWQkpL2lELX7/VzdEMKHqPuHolNvPeeolvFB3NQi9swzj/yxwWT4HbN
96JXYvfOgYh9Sq8hYy0ZLTlWhNVNfb84yhB90Uc0q8bzfgYCAWkqC8FZXXSTjzNMt0x6Qxp6a2Ez
Fr56p6IponzYnNOifZ/P1ZMVirMhWIr1BVjNiiq4Ge+fP6FFb5DnxGtpuQcmyGyu294H0+3slSAz
CcHKWMFCgYz6AEiYQBqneHX02A8XjKTuqHqtK2Fksz9QQ+9cy3kiPSAXM7lCLgiPVQZafxR+07ty
yd7ZOQ1y6FUWjym60UZHOchdyHHegjpAOkMiEkgBow8IHDW0LL9er/J/E/ZW0UjN9iJq6Sis8NIP
NnY9XIQjLtXAi8oFKtRTYz0TsW8ewU8QuLwqYH6KRwiI7mZgX44uiQmdQl0x2EWNvtGQYvKTxu7F
776Cs3LOYRqikz1PQJ3HrzWGTVkGb4JPPWZYM0Hyyoy29Lpv8qCXcLc/I18GOBTOeBCSHfR5aoNE
ibfSmSziMqaP+mrVAdexqm2xe9wGkBZ2Szl160Ex9TU0FKDbU/rfiQYzcB82HJMgpNQ/IXAN4b71
cOr5RL46LGM2KJIqh7BO0d3LlBTtWv4Q0b2QNMCvUnIugq7BciiboAjCZ5zniggUPjlD/E5GRc9Z
/M5TwMJGrEEbz5zvVfZSFstk7KkWW5AxXoSLeS+10LMoaGyN8LAtX85llxgY8JtQeaQ3svBv8BLK
geyOPvW57Ez+TYI55N6u7jW1QJRDuQrw5JV9bjFnYd5uXkaH4eK3Nq3vmFTGwLvnOJr9yEKc7/O4
PFM60tVf6Lqg8oWsx6bXq2AZMQsQBEx+b4H3dRHtt2wL8DOw41g8jKyN3LTQxljLnnvND8NYl+nQ
JY+cv8T8PcThWUsPIAJSPBS3MiL8asN2sTSfRMIKB+S0Db+ZVLeb4l/0senPRCgDoIuD2aIXmTjo
wem3PDqVfWORCPIyQxJryG7VohDq0N0l5KMZTL/l7zb5ZaPBBdHc6Vqfcji7tuZPMbcC+5K3enxs
5ZfYvnK24hLw0SLml5nZQq/Qft+oLau+xPHq8NAuYAFJLUfFD94bmLIBkdtdqnyXLz9me0+Y0KCV
bBPVHMFbqs6TEUoT08ITgIFkGTnCnT7OiF1zN4Z4b5RYzcItDNQMxutHmHips33hkOJykMyHdUyi
bKhAfKj89wIsWq3o92v2/1Xkvv9+O+erdtUfhoMMENqqGN2GrabIfJoV3A5/6FQSUT1zHt1v8IYs
wlTqUyukpEriGKY15K6HnaiH9KvkxeDrL1uA8xUT7PpLJNfWe1Tqgb8C/a+/hENEXY2grU25ZkYL
I1GEfBRFeisbe+tSqJsq9XMJVAvd09Qgj4KxZp6hgUm9u39YGChKNnHNfpYuY6TjFKCHr56RuheP
NUsD69uiW+vWdYWmAodduDwcRBHREjSNBHGhIHyq8+fxkyQRTvY9KecdOtRh3ANqSxH7edfJlQeJ
4UMpTcEq3HmqjGAdh63i+6I1X+eAl6dlHxI+O261w+zlHlUxglLq9r0hv0HumYpagNeGIC9KgOea
O+ISXe48Ps0MV4cDsrDT9/WUy0qN5mRn5GQRwWIbBBYjmAPUAynX8exPe1WIh5QyzZJaRtXL9sF4
W+QeRqhuxExw86FNSmWOCJrUTNYrkF+5ECtLgTcyBx0dZa9Lxjw3WeX/i44z1EExBLsq4TIvXxV3
BTPBA7DFijJ6H1/LKAzFuPv6S1RjCatkFEvvGvKqmZu1TtR6h0X16t8uOa21TNtybQyjfkr5NgrA
k3XzAOXLDgJg9mQ6TcG4oh86QQQZVXhvA+9ntcaoGMiAzu+rR3xuP/6OwhyJVSIijU0EypNqt5VX
kaOmxbEt3iKS3I4ZSQdAiBLO3CRkP2A7ItzUwPJ5cpRa3hkx+PVbHOJqk1AdH0FChWyswoeG2CTE
No7rhML+vg6o/zdAnv1XzkZwubm+xbLeu8UCYFOfh191EP7JMA+37D2/1HaBjGTHj6xLtkxlvq3B
BBchl8/8AGVucdNRwZjY08tCck7CJhNONw4+QOb2QQjdDaCVrj0H4R+/CxR8HRuK6OfwjxHRgJPr
GfTI25f0UpGioMD9B8rOA79DLpHwpMVo3lMWi11JvgY3SQDjvGnv5dkkrXkafgpgSq/4DtSJCOER
fXiD81f/PkxGNOrzvdr0Us6V0f3+Cx3/Ajypx3v7AweW6RQgvKeGHCmeSZHkMYvZkJq16zih8c6N
9fYhIgAK9WtbkcKoRHG2UPFSSGL2yXL0MQMd/k1XEhXJubv/6c6BOU24p4db7iHA9FLkubyPoKF3
37VHnmv95I5K2LS9p22tckmt4CI0wisxmDOJD1cDOlYs7cY7CPuY32IYP7L5B7yYQ61GW9bxlx4n
stDH8b/Fqh0FOQ/uNRHg7WmZ2FZZCSp5H5moerM8vmnCh3/dJL0LG7XLtggXsyFyEwUYLqN6xI/7
f1czYpwZcjybB4MZwyLA1chZ2PKaVX/MYh7spA0eQsrZsenzwTZjVurFlVDgyvRVU35QI7WiVxWJ
Z+s4i2qnsZliRxiubeo5GsiyKeQqnF3tgKfauN/CWJP4oOJT/0ki//N5hOM/Dcqt1M6+iIFQVBAP
OQHo/YwMPGh5S/krxQhmgTbR4m5KHo6/So/bnVVCg1+oOS89symJbkxsORO7IcKW38zE246BwZo2
UlqdoIoeoLYkY9AiDBCJoq+7S2iXs/f+WEcPHl59b2Ohk2PM+HELT1F852lBzcbaSSohhVa/leiy
RsCTsSNF7Nxzy+9khSpBszZ8/5tFw0bwWXEzu/quKv/wV6F0eiVuEpwx5d0R+8w0SllUg6cyiU1v
y3XJbecGKBrHs1HH67eTMGMagAgpalejs8w7OQPMv3hUjTnY41YD0oUxieSn2k4/pT+Ex0EUTAID
yYaZAkifixRbQjdpBtiNJtwdh3VtWdXzmR6vS2m14COVVy9gkc3nQFBLtPbj8wjryzFpdsW7GWQ1
0ItUrbk1YfgCtmAAakHOPtFtXHDpiODltK/8WXTd+QuGqPHJKhvPKHpxrVEiDFacytEpe8St2T8j
sMwMA8ciY6AzLF+as8quUlREeSUxB38Gk1Vm7JdiwKKf8EQ2UTjAzoT6Ig3xJutt48TGFQ0lzmp2
VY8qYQmvYSKfwaykxRC1uviJe3jyLwDnm8bfSzEuuHNyEDZqa5GOZHaF/iiEdwXgOQeWZCdAK6SM
K8/DMtL7PuG4rPZ2jw4BZUnzU1OqXwL9o66Ecdhe7fGpByhajnsyyJXyMtNlvdO1zK1mUd3v7JWX
qb1R0rXBSCrYDRFJCQUEIczjc6eoA0jX8z3lIvPVPr7UR+oIqPC5JUa4OkxTxOaTU8j3V1WEGOEs
r/gNY12W03LnxHavGng9MmQI/PddyeOsSRB4wylndegwgR2uEv9XWKpEKkK9vn/a6jUH4OUKo5XU
dYpYSmVMHqMAGTKAdOxXX3IBIdkRKUiEDAK0Q0Jp+Yun1J75QQ87zgLfkoaFamKwJU+5q+C1k9mv
Rg5o9rvRSQ/opiBfN3cPiVPZniYKmE/l4lXpSs9knfOaj2Qdlf8qrRMVoiY37Pg0dC7IlOjSgU3b
HgBsNokqm42HVLYM3PW+Cj7nGms21xVxM6ScWPDcv+1DF5D5BCTg5Kvmxk1EiUgBXrgzaIHz8VzK
eMeNj15RN9Gw5fycIM6qbo+blIWk7Q/OKxZyrt88xmqw1HdmVjZDBqKztsuFRmMnUFbtz3EO72An
g/mYrq75g4Kc097i4T4FOeGzNpA6rztmlTSFZaDvN7miUG8IJEWvSQMczjE86lftE5Xd7LR+8tKv
zdGUvmCVcVyVF8cbJiMEmglZd3+YOXyoZ/0VwgOL2vgXz/s1dae4/nsYPlg6QYxPU8asBNmUk4BO
HOzs0trh9tqb2Q8tosTU+FpVO9h53DilE79tZA/ndS20UTBxu840B7X73077fonLwFEwE3bEcgA2
GIFbOaC8wdqwptQn87+vrlLCfBupetYoBacl/1OnBywnNe/V+MGnGqDywVu12sJwOQCr8Gygel0l
1GgLz45SZZGUFJe5ld94+2XHnGYSZXGZkVOlUhdk39Iy5pdXrqj/fMx1xCBdSvKGclht9FN7T6ac
/E1bijMNC+zXT94I4tzu01RDNfiNg39lQAtzd0Scz3aEXyWElanTUfh/8bLvd98sFt1KZ0WthNKo
GWYQCidevuOjPslMGKGSsqD3QulGFqvbQ2O1KGKz6QWDvwlFZnhFYfDzXuxw0MMlR5zSZGjCzo+p
PuMpxB132I76fI1HPs+J4x/VU4fwbVLiejsNw05DYg3zPqBz/Fzv1XvSkUWj2I0a2WSyEinwQxFs
Lle8yoaIIMjfYyzeavdeBh1Vv8WRtahRp2MiTCnD8ftI3Wi73M6ltLcFCe8nShP9VQVgWOGFDbqa
GrJ3A2qa1pJjaQPvbxECVNF1QzHNY7NcAn2ppPAxU3OxuO7ZBWFGR1wGj3CAj936LKd3Nc0mPGJC
DzErV6BEu8xHzZJ0aaanaPSseGJf8jeADposNR6Xi05paxnzV5R/QM6MwB5FOZCPZ5uxPGj75LH7
bl1BZHbqM2rkLjdIm6sBg2JevFGNL1hAE5UUumG6c2CAvEhTzLrK7D/LHbtxDTGDKxqdW2QyZVo5
k/PO52pSgtp/Qm5/h8CFU6xL718JPUGuuN0WQ9ZBPhtoNkJqiSqI1/webnogI1Fbzypaw0LpJld/
rzqfkm3+15FsA15yZRy3G6JSXt+bsfgaCJQEWxx85aqv4rAnx22lQjYIAhd61sqmWCMrgFlp1NLF
5H8+XdTo2+cNc3NwkpBV+eq4ZHlos8AYA+iEBt1y7X/TwEbbPc5Xnzt0dg3SoL0GV0BnDB8kAPBa
pce/RFT7Y2wquTgDmxEevdEgaRxW82jWu2ly3E+lv/lQoAjclT4kzg51UHUWA1zZa7h03G6HC5JG
ceyVvKJEOG3cSu++X+gXJvEaIWWXsx85cbR4jLuHFCz/Ff+Ehdcxt6edL/kUTwjk9gu5iLYHBPOj
2Ge2Sx9ifc4KgEEeXVNS1ewex6xIWE8z/+Jt5G9WyfQDl3iA52zx/wfH18yh2kDIHoXoq9M0+83a
JugaTCDS1h2UGiEFBbReXyfyHhznxE/L9bbuaZh7dijt4lJzeCYjCkmDQ9VgBAwpxQixrJPYNlJO
C5Cr/xrF9DqXKfYAmD8NgUvY5EzEu450hdua3/iDKMe4lLJEINQIscC/MRp0flj9JIHvvrzfA8XB
X9UOcRjIrtPgy8DfOq6++oGg9A4CnZxcofAMPgnHiJfUmLtIafiA3LAumrB1y+ctqZnTllvHyuwZ
i+I20hGARge9MGVHpSoN09yqlWwdfgBXfv9nSZ2nSL8VAAOwdmz956rhU6mtxGQkDPQ7aJ/FCxXZ
+3RpN7efYyMJflCg0nI4ov8ZrJupW3vNIQ+Sl4xxD4B8l2s2fLSr6DMlHdPq6ZCqNcTywDLskEKC
FQYlFJbM+VK5dZEchmw2Rn8s4sVxteGRMMkO7VMy02BbtpScZTJpJwgl0RS+s9g2ZErMMDY//f9e
zErJfV8VUPaFq25q1x3uLWYt7XAO7hWptUTQfAvkyCn9D1MJw44Wfhq/IsZDoxHcWFvMCEqjtkK+
kR9djfz5B2y5tYSFPwI0pC6dyUqVChKrN5YsDqdagGc52KSyJQPb1xkxzKETMQkGN7BdIJda5Iqb
xDP0VMqxzTNwqBqEcnoRTqU7Cp/zPMHH2NEtq42NJ90rhNOy8qbIWC6+2mT0iXKCJceHfOnFt3cB
O/Szc5kRZzJjNedYzv/qd/YTMBus5Mv5oMbrWUF1W7CMHLgfqtwyed0PtFCGJP/Q/uezI2z9XJ1w
+YKUS2q8w3UClVrGSYy7I2MLioVHTTn4WsfN4UlTNh/wN2XGXd/plwNZ194wqIvP8dtP+lRoAG3e
PfHZoXKK1RxVOgEe1YcPv5SpO4aKRb4eEQqtLYBuKFL0RpDqtmKnH9lHv7SbfidgSYFTneY9YmMv
nlR6oTPuZCe+MjTSus0RTlMMZt5y4uNi69xda6GB1C5BCsPe9Ie59Ab7ouFsjpxOqSufH1YM7Y0O
v95fNHE7ecxSmmg6mvlBcwPwzpsVuVbgZq17a+8PI2u9oRyODhhCezdGBNKfkOUO2uKgprBIzl3B
f0bbvQN1+F1Pd3HXOeXTXeUchSlEuP3Cbe47G1TgA/xEeAd7Ua3reglmFdCkWXry5ey9QTKFGLnE
yEiLHy7KEaWdB/MC39mvXDOkA8WAkle/WwfyB24dYArcpq+oOz4j4yRXqrATlHlWtEjNrRKvx6er
bN3CU2SGnUgRkf5s2FTf4eer5o5UCJb+hgqn28E7eX78QMycCM6Tixe+wAIMlFjrvaWgpea25WUa
uG5znisAKqSaXshaaQYJjmavEtxqqrq6eIR1Nuu2Z8J+a+yIqWTqjvg1QpuegLnExwCBYMTwRb4T
J0V92WWkOB+D9ovQgsLGdLJjV3QH4z71wjaNsf5wi3rd6tX8rrOIyVbRg1ys2ktMgalp5Pj6CQ5t
XYHfc0DYgZn9euHNGB6+PYhxFCxcjAlQbXjboAr+fJKX6gaXE/vjK5zKLPqsQZ/EFsUel+D63od4
YlplNVynZnGy4YngNfyRlm53W7fN9cnaRMEYBSDcCu52W0ECKiujghwFjIfQR3FENOi3Hd8WisGH
qGL3dRR04qNy8npHoF9/luvWMlVhRUPxG4POTJQkGRoQRFgPO9BH73wkGHJ9wNRyTXSmkEWDx6an
BcCz3AFKNYUKiVP/XDGrCVxi2evaI+zO+8te9am0G6vNXV8MWwiH3V7V8H71KMlxbz2as2zT37A9
kkKTvlazV4gmLzycjQgF8I73bY+Xi6J6XEu6kLgCc19f57d1ffal78zHSltBy9TrM5Mp7kSf66pl
1Y7HeOQ5bL4Qwtrf6HA2tAWayPQPRL9fWqxXkm+IpBqenghq7MOP2mfZ4iqAoqCuZwJyoOU/mo1b
Mx8s1T8LiUTF32KziQm/Xmvg1p78WIVOEUujPILvGte8X2/rA8xwUU9Ent7VzlyM1cEEzL08ZEpL
PWvVcvHrlDKZfbWHhT3GcedSrUpDmSq6qft7GBD7Hj33HvCMOs7F/xOBpKL2ESlklkTSoP/ECB7P
KaHcF+p7AtW4WCpaL37jOV0L6F3GAeaqB4kA12/HktGgPm9CgHdl57dGU9WscrU7i/jUa2P9Y5o1
kvX0Ey4RM5YBHBPNiBZ/JjSddcDmfyH1GxxUTfR5b0PaZVqZlvrrd0l6tkAPmbNPmr2irIvG0BEM
7THcVn9Nn+jel8H5xOjfVZlVfo1y453YQW3xpSFV1VC7HZXQfJFTdGk7ihqaluXHxdELndttdCZI
BFK5p1JHJG7vGDxRUdp3pBL1jT6M6PqvOQgZMsLI2MwJ1x9NhILwzjjU1DbmI2VTpr4eMiMFHYhz
GwRPFON9XL43ifXXi74TEw50gJtQ3v9So5WTr1Df6+jMbS4XIiIL6XBKKDXBTo3d3FJpqVt8kZ6A
kSeBotlkhIzFA2MMjB5mpFCF/lOyS75x34vT2xIxzH0jRXe+hQj39IMen10NDYaRmVDbdtoa8iHT
gRz2pBp75RRpcPFn7+arWju9Y30uAniAmRl7+U5tIROQ3/tnbONKqKeCRjJw1aYKU6I3c/96ZFFn
tmAdO/0J+nfjDZebC/v5Bi9Y3LfA/KlCedAS8Cid4ahzjAVB39IMrGPWm6w6lbQZQdl7Us725kQC
DQbkf363Zland2wJdlbiIcUaNcHldU5V9lJdZcnKxSB7t+AmjKcRbrLxEK0jhS+OtiUhotZdacDv
S46z47nu+/5YktmP95oB8EEVrh7+DQtDt/37XTQ5X3aESIGspJQ2H0N2JJwHdhrzl9ulxH/jSkiV
ejWCveNfWVSL6CpRzQqzhyWz9Oi/79GFmWH3y23UCD458+t9B/OnChJuLgbxoYof0kvSMmLJYDIT
vLTSpAdA6DoP5/fwjLUrK/jZCviWj7mUf48sut2vNWl0KX9TWAWVyfSe71s5fk7+V2iLTRUsI37G
x+kJ0XMbuiyDLLyaSS1n5nqaM6cN4/YnxMf4K84AFj4hU5Svzt61tvHVt2dF7iDPSCBnyQ91qTqO
AkRVGN3dwSReBSU6KEm/O3zmdg0Qw3lY5WxBib33/OpXUu6QOElj/GuyjpVAPEzxOQ1+9Ay1VKNw
npFzTQnSe0w57/+SXE8I2XOKK9wioboSoNoG5c122NrtEPlbZUf5/Qog3QWpDflsqMUw1cm1Chf1
6NVIILNC1L1btDMQn5TqgFfgTDoK6Eay7JcucmJMiy+gP2aiTa31c25S3dQP34DWkSMGKw1v9j4T
RMhwZQEdX0b6LrQDOcwHanrj2btY4RKrwVniJJhJIZowdYi7uNtAuw2oXRcP6aGP6BADBqJ2gRy/
qMcVvlgyWP2uW72fHxhDYgYBMFe99BBTw3XlF3tfgS9Du4dkIG5qe1ySMiRIs4gCYLZ5kZOi4QJN
LRFqCyBmOqtlQTzw7MfrvnsXHXF/Nw/BlpIHEyZ8vOlyJDMhvMOlY6vi/tmj/7xQqYpsn/Mc2zUE
jxaDxMgLYq6G52PPDmGVKS1xaYFPKwpuDVa4J+3TEOuy7XrdsdBT3VHin+Xomq4YTestjd0LImaW
VKYg8EqPncAqTpy1lvB1Ej7tHs5QJ2c6zMTF7NPJFqAMQroS81DmNk7o457LPuo/UBck6PKRR85f
1HwwiY0YSA2FRBYRiTJIwT+DBlCu09V912HNzbUmdRHw/EoGigfsc/5pBcqxdU+g5GJERChY3IJZ
LV1ygglghBHb/yVPV5Uowhu+0M46CstqRGnRrNG8DnZFSV3MFmZTMZW1qiLkkXpipV26vO73Rqk+
UYoO/iAorsNJsbg4vFHmD5ChTDbnSyopW7m5dLi65OiLo7SIx5MB63mHrmhgrBYFD88SW16rDEkM
LRoicQuKK1i92TwLIoV4h+ZMuIiboSGjVGeXs7cfBPTCaSrNeP3fQd0u/AuPMN0gbsDs3NYQhwwO
1l1uguoopc/gXsQGlA/W5ewBHPlayjTmAzIYcHIAQvOoXoc484c/yUI/P2y+rdh9zkkpZonQxDXN
BkX+WKsCI9V2FB+vUV3lbuiKmlQNz9tUEZiwrGcKH1mk8GK33iIv6WjwfkUmmw70Mkq+k//3/iUY
RmQgln+qhRhKNrNraUEOE4+Vk83hkjiSgCzuJGcNpx1bxKhC0YAf7ZK6WmwGRpZHDNBUZLiqnfVQ
jPehfwOK7ADDT/liWaqyMYzEGCd0nR4Dj3DsfOeiQCZ7qHAXpJ0Boojxz22IuX3qfAEJIITVyXMh
0QA/iJsSyuSDiSPX7HKgP0P1lXizx9PH76R6OVkKr/tNYYNwazxbf98nJiRnTFWFDnUZw0ulR/+D
RmtliP3l+fNiKAraXoq1XtKE7xfDsUNxVBsiT9nj7ZD8MtaFGOq3S2qFUTHQnm73syS0H2h33JWC
hXgK33Be9ehTWojcvIvDyMAtz/BkCmRF9TI9VXKNP4Lz6/xZRtcbQxbojnophGmreAU9Ej/MZvzM
lgCUr+rH+NwSjAXNQFPlfT6RVQpGbQmSH50rkY/SEHtu/FrwrkBn/Y3QNgs4fXktlPMqo8uVAhKK
+fhZY5DMZHu3ewaHNYtavr6k/wB0dPZea9mfiJRcI11qmVpD0Zl+n3yugL0RpUTQFdr+nEohFLgK
PNLB9wbX1QR9OkSVoPKWcakLCQfGtLx7cSzKqKyweAZ/+MUjTIoX4DjtGZbeavzA6B2c8mxpjccP
T1vuSldQ1dheIObCde9OdRNVKvDCtEabdpHRH32beTQD2cGwJ0JNGC+/UxhwDYhzCKgcYgO0/2mI
KyGH2R2n3uADemI227xEbYRzP1uV2lr2jFTkSjrn1NFnmfm/J/jvEXGlEJZP+mu5teqUnIT8jnzU
a2s5EAnfUmLBAnBW5Gta2QiOy3PwLS+UrZjeqn80uLhoi7d47FeQKxXzqwAH9QCZ8KrGDsxlRYMe
mFoQocD/qJ0TTiNB1BDIW6CA7tmQn8NiqczyIwfE60T92Y8u40W684dY68FOARPcx5/M3Qs51yz8
p9Nllq8t26kRBKWY1mexHgLY8TcAXzUILOmg637WyJi+JXcL4z3ju4dX2lsXZHPeoWIe0jaJG5tW
rwBCZ3k9YWLRR+U0hjIpw7unpefdg5ieMsw1j2u1edKz90zNAs1H+GOyWGe9j4acrcnDOpxW6FxY
bzlCZMYxdYZEDnio79jVwBzQxhKLq9jhCeBMh0R85zInYBgnM5ITMNB+TwF3nbz0w1GMc3D6bttK
YNi9qGCxMrHzivl8sAFN0aLyXPS5pIHP2ygFtOTttFKuWcShTCfVPZ9ygU9nb9SaMgfgRvhjPS9w
PRfQhMeHGToM+w3mDS1JLQ4wx+UX57o4HX4oJLlhBn3JitHNYRX14oTGH/8uFwcEw4Qx/zqzHbGs
K3gpA2ZCpaZkyykcFOMquV5ojBJOeJayjpn3oM+qqjq5Bk6ALU6iuMtD5z06qPLqdA8HiJ6PHY1I
XwdNNN7/2om4naQ8qXqk2jSnthur/lnF1XIt9wwLtEN56uzCF9pVcUxz2CaHvxgNcX3oNJjjy5QY
YM+5vIDDIXJ9e+iML19m86vY2h9ZOZU1Fb3lf5yeWR1dspr0MiGH2skiMNzHmvW6wG+aO58783tt
OwtT1MbisCs01T5p5Ji0q3RF0wf9YsGhhj+z62GDlz+Vx5+uKuQ9tcfLQPI7fYfNxjHvmAuvZ2Yr
J45RuNsm0r7hwKr5NILaQMcTeISup2ZAorlTGr3MdT2hajzj8/jBWOHbVXeDT5yEcXVTh7x88TZr
+Dw903vzIOu0YYMWDUAVsBqAsdEk7cHet/UvCjl4CfR1OcSlt83/kpO34TytdVeQHFJ8jAt2JiRd
hzCsW55vgVfzGDIeZUNU7U59keuvbi56RKQOMWa+LWFkdZZDy8LRpI1ikkkjOtslpnHQtgvcBkUd
hpyI+8cLbkMRoGGGNW2zRsW2WLIvNR7kKjDJZaurP2D/M8uW62C/f6E2W/CV0LbBDE/7qq/wNjrV
0syYNPacludNPyigVgJbcxlUNv6sz1KEFgRN42+Vsod/ag6VjSfpLsMksjbscqRIlwEMSVBPlFeT
ob7VBc7LoJf6s1KXxD5BumIK5h0E13eT5duE0nugGY/YMzmyOWqwfZWb2pqPXSLCa9FLCqWzIFiX
c4U/Qe5yp4y+w/eq/fqSxOX2TFacFw4dOxRc6n2/pKjS7Y7X/PWENetT3F1afeCBlmrXBAA9dGGb
ZisdMz5NRqivqc4XA0xmU/+JpX3iwHYCHnR7aqU5JF69vlxeYowQxfOZwjC1vq6ugmBwuKwnk4wy
QSRhBVM9P1a6c71Gf7sHQco6GnK9LFpl1Lh8wp4T9BQcwZWTg84k3gU1lksGCRhVi0XuGL3LeStF
V8GShDQEackOtQaKfVFyejhmnqHbNLG6+pRDgFoRM/KRUfg4wjrG0ih3VcuIJi9tly3WP0648nWV
QOKb30xuC9JKdysoFNCKkFzAF+DHZ6JUPhWDBfIZo96TrLAQjLPUgjfFoq5dm7amITjZhYBZ+cuV
vXBvYmwhhS9IPB0dW2GLf9VI3e3gOBZt5vtfpq3mvbZlMjf/XGpp7g7aRc6CbFAotFlgBvhc/J6K
VHj1zeZFqmoWFRqoidRzx9f6342KoAgw0MiyCuNMJu0RUoROJKbAthfKI1aS8/yXSKxUjkIHr8nk
bhODieguxpSuK4KeVU/KZ+p2zgSnhNSBtqhKI7WM41yKn2rRvsr9ck8fADAX+Fmg/hZYPLm8Q2Qg
jnqTEjUxxnjK5Ldw84QGNEsbAhX3jOjL16fd/M4LrPA9JNoWJ+p2bVe/97vQzNfpIe47scgPNOVY
o3H5ov3Z26P1jmRPSt61POfcelEmPgvEi9ZrqzpIfLOYktMg9KjEu5KcmBSo/R5dJETDM+F6PTsf
LDFM4aFGQo/yW2PJla/nTc7rR5wuFrU7EGtK+MiCttiVGHOH0qB/BS8o4Azko0uVf9UBKz1Nh0ek
gJm9Hyw8cBDuk8slsgKpIhpwaHNIsaOr580ySObbbcU+2tVzBJ1HnLHQAzrpKK82HKErVPU3uW24
X/GQFmyrAQ6aG3sijTWT38s6oJVorOIh1jwlSdtoddjV0DaNBl0BHxkI4iHlJtCZMaqdGSk7wLRd
awTgnj/xoZAo9cOIL2XVPLlNh1wOZI20KQQpf4CXYBxLPbv2K3CEB/JNwHf22n1C9y1OKhJLDngr
s8fEdlmG9cgO3yGcOJD32eDmfa0MOBijHKpWoCXO5IvXtW8FpvxqyMlIUwmJgrSvt6fsGWGKbbu5
E0Xm1zXZOMEDFuTlRrvGuPBoy1oGDPfFH7A9H9Cc+BXNMzEMBV36FNc0DnAU9MpTkFN6Tr6/ZOc1
RKPCn+0UUBSWSECsRnR62KCLB3LbA3X3xcqQS6ladBryVL6C/N5ZhkQMH2dtY98+o3Al0X8MX6sG
LNSs4YZaAqszxTcwIOKCNZ2unieMH6bfGZhL0h6zP6OIXu7zcyTS50COjZP/37p7id3MOUX8OVvq
m87RHqZmCTDlpzZ+ZefzKQ+x3y0dUCAtzYzrc+VV1kitcvEH08OHLnzLJaD+JVZNOf3ZwIOb1Am3
OR27Dv2gUVbKqBK1tXta4uc39MjRDK57HutR20tUcT6L/Sg6ScINSwTu+iocTMFGPrX22wtUBvQJ
zEsevaKVD2d0TrMHmmp++tFofgIUzqn5kJw7o+CCAu+TSx18nzyf7hnUVM344dHTM2d962/OhxR5
+Q115ZtJbqDJgMLLz3qexan7ev8g9IHTHCGxM4HhdHjeuDbHBi7/XK/8S+q6/qpBZoBXsuKPgGAQ
DI1BC4cpFLiA+BJYDU83FnIGUEI2Wb4klZlvjOGv0XHKvC0FXnolI1krRrkR1mkK5G7IM+z+oIUl
kFz0cJv6F/h2VsXERUD7MaA3i+t95mC/ThgMdGrFYn7p02g2JSTYXZN0ydPog42zq46sElCSywbQ
5XZrqdXzN8/pbww8A/hs4TF1gNlJqVuboJRYZo0lOZYHBJB4smi4Qj5TStRrhFTwzfIQ3FrB3/ru
9l8E/f0P67YzxUV7ewuTOM2+5SN5M5/BHVBcKI2MINHKL8Vl21zE90LSZl+3wRGmORP01ngbIDyx
J0BFDaieAIKQmsf3ObqP8sAsg3bf7DIv66mdVNFH61cJIPFfi8G783CZymtN5UGlWvTcJGn6/lSH
lzwa2NbvoMqp+adDdP6x5NefijBkkI3yFobqdUUx4997Qgn2Rac7pEDaSx6i+t8LigQAuuS3PrW3
ItZnZr2b06RUntDkmpK6Wnz2riWE3L5oZuTssiZpTb6ii6LUMoKZ3tH8EDfRpyiDz/N3JaN95JiR
B7vC4SplWIjis7+6bKoJ3LwKpetRfYdQwojAK+qLYc5gAaxxpFpK6X0/uRPzFUIZMdrfHBg9YJPJ
hKDl/dnPkR+KM7bGwe5B+vbPvlgABWUZeuG0eGy+aPZc/ZeiZCwLsLpqQbpX9fXEnhoGpU8nr074
b9xRUzwkW8HvWRTbHlwxskPqbZWEIxvJDQC6UYkWRRvT9pGT0YZKPySYjhBwqOqhILixjuAsrRaq
5eYXudlnWF+PrzoxapXU8HgXB9eCAD+POSJheSFijd2TyHxkNVoDti2d6KUE1UKW3c25TucHM8YM
ZF2/9YeFMGTNWXP1fdN4a7fI0HSSZ32Fy8iDYYyJYEzx/5jmkg4y+culvgpJIhXIyVzb9/Zznq5/
/m5Ir6NMkSLGKyUz/ijZoBtKX4KoWu/c+5M+xS9GrzmRaBB+INpHpMZAPVDgdJiRiNvXvy5zuson
8aSfAUTrjBxspp43Ex+S22wEl+7qRQy4CIjMrZBCr8fosZf9trazKGN7o4eRXJALo8/vHCxzhr9t
RRGNwvk6hsNJ1IFjJGVuQtSzqP7eKgWzR65KSdmEn98UyiIJ/wnBmbHZuyR3XLKO4/fZC393Oflf
vBStmZB1t/QGGelzYVlaDoHHAeqfhTBz4UjtvIqe+jf7Dgm9MKilRUogC/ubwUg5edvU7m2wFYvC
KwXDYcf3AuGNCPhYC710SLFEkPpcLqbUToCLPPRQEXRtPSk63WK53jGKLkytLeMzuhcg29yJz6Hl
reMg45/bJVtg54kRbOdqnbK3gpxsWGcyP+cXpZ125It1BFZouBF/Saq9Di0aEdUzmENzxDn9WaQL
OJcwW6sM387bIhw7vF3m1U1ByQLc/igh2l8dyTnNst5eBYnmXKeS5SjLhta/kio9hH/r/kYVKHEg
z32GuPqa0Bt+mb21FZPAxeLNu/rEuJKQYzjNXq3gPI+bstdRb5E5BqnEyTqLXOR04F34Aws/HwgF
wYGy9THbDYqg+BEwoAqvrlDaiUmd8xg5Uj/tBr6lBxOwUxQ2e2j8GAFPuLgbnhQ3NXW37fMdoP7a
7UXvIvldrdQMT5OJUfXE+PpBD8lFDW1Hl1sFBd6bkoPxsFkKeDwIW8uUAhZa8C1bKFTZZn0xFJp/
qA+wSqxjMwBk+nKfEVbAZuaLKKeKMcfNQU3d8rnYkaufJLsAg8BZXwT2x0Waee/0mahrFn/4fhvM
7aCrMo81vqzoZ/1aqZuaCe22ylMRiSXjGK8gYzjtSR6Rkc6O5Vxv0rIvul0Hxo95aeaomgLW7GkA
aC2sx3yhIVHHqf25p+e6MZmBCQXaAjx69iJYlhHD6Haojm31KCmSDfrMufySoVckdMIUsc5V7bPZ
sbuDJfPAx0fVMRXoT90u9hBUddx7QOvHgn+IbngVCaXH58+kAWNPjzPRDGZ5Gqa63cKUwID2UyAj
X4XfO8AHThZk1D/Tk6pgm9hcBKInFSVRs4iCp81AF4rnqQvbAYthsAB/tW6T9H0kKRMVo7+ZjBFj
OGQO7t75Q1OCQS+msPRc86yMdBF3A3ZPc1vuokJEMJYuKMsYeJL188VGDekLEXRo79CcRO8Vnbc/
FDbtwra9Z402/WWv/9sG2DoPQnizRCdI1N5CdXe81yfyh7aqt+vAH/Rk0TWk4IIiiejSbY4nYlWe
doB2uuIlY9gJeiIDeEF+PeDHf57J9RPRZbNMOik3l/dAQVpxxTBsskGYgbVG2Iu4r4OTLFecjk28
sG/z8natU/IKlSPJHmF4MKEbe2d5Bpvit7K5KGZ5ocnmc0NgB6qzyXi21Y3Wqy53SFXuPlEtnR03
+5b8yOaF+fI2JkZqEfPddvMLIgC4niVcVKxv7AgELs8xt3OFEgB/IMp9awhxiC0XkK94HmfD5T8r
s+FZwY9EZL+kcWf8d4DNCc/A6TDWgSgEcMb0nD5T3UWjvwShyGK4l+lnyi76zq5yp7hHuSSK7mQT
OVlyGiWBoLervte9nwkchAjQq6+N0vIZxx3Rsn7s61mUDB3cXALr1JFjv3qmXh1YcHPSUkpll12H
k5w/kmLmIeR+8+JwuHSZApgnftrdjPyLPub0dFxHlsiDAzdEbTDwqH4WghdSTg1k6GsQX2lY8yoB
GAnw0wQ0bJumL03twf6DwEgL8fmy/wwG1ILSf3GXKFEW/rBfvIGrkn55aEfYpoQUcTeCBrwoWXOZ
7s3l+xnxxZAuMMNrZp0kjYHw/MznD3oLKWf2yB3cvNOMvRQoIXLp4TXeQOrdyitauOrUsmaoHrIQ
3+CjU+RDZRIzkxui6UtIP6FHOgW0XeSHngdAFtwkKf7NY8K2PJWDyv+p3Na378qCTxjepdZUCzRX
5RKoKxj3fKOXc1AziFAILHhgI76qYgBWVWOy1xpF1Tcy2bSGdSnPiwzddp+fzR6/mdizXEnYPc0G
Iw1q7Kd10ljO0pH83c9iSnIezsDV9bW0Nj7SlyE8iM1aRNP3lNoRlgIc5ldRIBI/Ml6f965XK3KD
kzXadaN7IUi6BQPLfh3dMSoj0cGFES+mMm+vVZnXS2biMII9Uno+JJrzpfFp+I9XD8FGX6JZfYwp
+8Rm+f4FLOjxzY9slA1JIZ86wYEX+vIuswwdN5ajehfnPOxLDTxWlB83Zzv3bErasWbnLoXr5RrQ
1OiZC/PSLyJ/Ro7ByNj3hDuZQ4eA5HXZPU/Az0xPxBTBqOLFkhiuIk2AuvfoofBe/mZMgjnIQz3c
qX0AValEn8OtrRrJaL7HPiqMo2G+W1vMpOmNgM4gO7uqU8DJFrYOMrTijKC4kzfDcQa2VtbYzzIf
SJG9O2RQslb8PqJ3uv2aejXdf0jEvlyhZZ7HTatHvSWWHbApUClgDZNaoIdEg3oQBkuZf6sz6/wO
YtFRDSNuvjyyng/cFt1o7YilBRShbCSzcnwVyOWI4sSrottWI7gQ2ag7+4nZOTIYe/DlHrxNNKx1
YX1AK+DB1z6oZb1iRB9dMGCaF0oDciwgnWqSgFnJtWxbV4lXNkEkfrNSoe/irIowbQlyVV19NnIR
b9ymgdgvMNhm5zJxK+Ni9hwWLSBxPD9zgTa8dnuCy1mMDxSQWfFhnLAVIVeFNraHlyZAbHvIrfV2
ZGMwnXbhGfW6CLWYSi26IKw2f0ZbZxd98KTu7+GTUi0TdG3PLHjwyGxYpoZEz0yXZlSkdxnfMXsa
ruozjtvNbpTaoywuq+omDfmRsbPY2MJCDB0OUMSI+pwDbwclk2dY0sC6TKDD4x5Q8I+8rRwv4c8Q
yiWqAXzA2hX70VQb+/sqdw1BdPo49Id28GLv2mEVIKYB4XczYlXAYr/O29adwwpAy6e2W2JSEpmt
2Cbi/gRfKTjxolle/gOxQUF201fOPwzIW1UtcQgAflAsS3CAHZOhxW/1yY9IKMYxWT/kXZ4jvdhW
QGGOwJOlluM9y0B+nRW+pO6EbKrT93LX+uh6tckUtwZbeb9dKaf7b6WtZ3+RCBVJrXz/+wI5KpZs
6xmb2jRP5KsjVkF/HAp22pcYvky0V706IL4QfNXMqhkCvU0ejIHiKfGf+cTDvraYrlq6Qf/5mpo3
YhMOxlQ1r52AKkW+ZoGNgf5bcRxF17d85XbcVX1bJhtZeqqtpCOy6UMbnBxAf38YQaautqjfXdKN
lAgtNz1URWrQ9MR906erCTsGJ8fH7A07WAut/usqtkZSbXyK1fLdIyFS0ITUXvOWoe7V2w3oXYga
fciUdWNJ98hYo2hH4WCsKyCggCDQU1nI9fqHx62ChRuBU8zL5252uX5nAofkyv46K0BnLaeWUT4I
KnjKIlIeSUzQ8L60W/Ry6DLNPrEn1QLEVPoTIR1yXK1OeeSV2SkGawRYJ2CFtaumLcoXIPDtiz7S
nOE2G6wPcQjDXL/tt0SJRuvBvd29ckXSWFfe1C30j08RZ+sd9PbdRaedFh/nM7Entaq9OAK8SEVc
yacWPWHDEC0YSawJq9mHzeniMRt4j0to7GSAzEPxae3agpuJBdSU9aug12uVvr6HqwjlR9dZ1VQP
fU76+DHICnyhYC1zVFpxbALCykKvUXbqwXQClrqET5Us13a7BOWzcgiws8Wtnbb07EPagjvSY4KQ
GQuFxIKATudbmRC00T2JaCwKqmLIcHMX7T8FXPIE0ga+72Fk7ngv3Xgb6ovihcxxYcci0W+T7do6
dGmH3Rfy9WbpVQOwaU+klUI8g6jbi0FkIjGHaeqIUePacRfvhqE4aomuLSdSr2V88f5MkBJQRXkN
m8JCbYIfEY2xrLUWx+Cnb+4zQ2E83TSemjJEpCH2iq6n8pn6cMtM4J3BXfQmhWwWH3F9ECj+pxZP
NbEw6LjkAMJiZL9O7qoz+V6yeejRduXXneEEyle5WRnjpg/p1+OsYhDJTNyiA6O3ukPoKyy8hUsS
3Nh5FhJ5YTSFTxieNK3ApFy4CvBvVK62Zwsn6BelkYJbTv780Uc6VZG4CmDs1Xu0ETGpUclJVQ8k
6VUyLOM3bKpPzh7pK48mr2eZJH11g5Ie1C3quC+4lAU0wfcHAtdyO+xSZgzdD0Yk8BB5g2r4MfQB
i7SNuaLPGu5v7uZdCO9gEDxfJVf+lxpeLsxRDz5fte3g/PgNLP0k6AgOT9q8o28AYXz1loNPQutN
xxcV+kjTjOoWjdGmE8ynSdWvwzRBafhSrRYdyZBZcc7MKjaUXj6y4w03VT8efIjVyglCx3xQwxoe
78sOAFWNBL/DlSBW+Y7oX6RuxMASECTSZnntdsvoTiiX78fko4zArJxSjx2OnpR3CNikHT6eXJjI
Q7ZL0RGmJaI+wLkLpVyy0hoQzHnlmy4HAThbpx4CzGBA6ahry5p2rO5mSSnMU/qRmNYOhHv4Z1DE
bUtBOfuVuxraEC+xZc2h31JiVA5228yQAxixw5wYwy2EMomoHlbtMOdbG940QJPk+UWQlX0/WAKe
VGcWyrptlTcGlrSoxjdiyf7CCJn1ffSkzH2bEkcpwMSYmu1v1lKSXrz598UZlHOyhRwp1GdzU1U8
YKkVtV3Qsi0UgAe8WAO48BIURXEk28gfT+L/c2gnl74xofqBLA2ADGpYdzos9l+GC+jCsfPj7eHs
6y+9tktTP5v5mIjnN3CSyEuS0OBm5Br/nrSpRg/1cK5y0bYFsVyO0fTILicb1HAcbvOc3gAH/l8g
4vws/xwBRQbTx7Y12ogxm1Kh7ZgEumbcCYwbJ4mF4SH1fb5O3LAuDhMuK1LwN5Ad7xgsQcq7yy2v
TDCrP26csrGYcZsiSM7aRA4LETjyvRhS/lFS3AQQl4+Vqv8dzBLvTOTfXenwackoftI4cXDzgU4x
AV9u8AfG6A6M9OW8v9k/hWe47lDmiUxmp+hR+g1xeXmEtCgA7Lx8N+jdyEEJe5uQuiB0O4CWjc5K
WI48rijTRLiwzT9JX3TaGYBmVlZp2kYPMlA/sh2FkUEtYr3Q4ZKZiWYcbw9HrpXLardRDT3expNA
W0XDInfviqo67LS8xRHKOdfLNeaXz0/xCOQJhYZDThLHNK39i5W0+eu1PuXWRuYoq0dbzy4Fv9ke
eZkYNba5fMa5FVVUllpbMDeKNvQTWgbj+jhtv9H/w1jT+/nIRJKUXtuXQBRP9e5N9pLeteF2445v
wknE7c/Dmh/bEIjuydeQONsqlwiB62riKCuSTefxT0Omfwml1pvaVkugJW854LWFtMop4Aa5IlWv
NRROFYMJw3HOh3IXC87pJwwjJU6kgit/9ZMmAF3+zLGK9IjrAu16A8/4Jniet0rKa/TXgYCWzJaL
za91L+WKiTu9jYJ2lw8S48VKdGU8iN52wbcfDAGdxby+5B7DpxPYAteSpEfSq/l3Vif/jvkHzeyp
/+wE0qtxmQsRD8wLKQwlF83b5jrB0HFv0x2ennymYSjQHcj5Ay8dBRPWd9rLxrfozt8xqPfUqjMP
2ppPZBDMTwCE2ZAyEXeWBQXxxjO/fKPEs7zWZxULGk4ke7IZwFtP6ePCfzrsnJ8CmHx7BqRVj3PH
qGmdHDcaOFvUGedJBnBjhBJ2HP5DHtyQsKRLhl8fddLl3rfzBhtuED31CPQkLdr8XtMDsDuY7CJI
InjLyel6DahlZ5Ow6kqFyj1Cv/dq7FDDCypYXu3+mSQhH8cbwq/xFfN3ygZNHw0h5xwiYgJdXMKs
eLEDeinYx8/koNMdfaOX5GaPGkOgrOfD3UkWdaEpYtYDFGiMo3HBQ1fE2UiXZpcf0shQ61cnFRf4
RzDi+awuqnWk0yg8vYPcOZsfXE/+buQpxTkEIbNer/Zm3KxWW0HXNPGCe6rNS0U1rTwOEmTMfxXH
JGxJfL5jV3tVQd/brNP5DXy9RZ4vg2bVN1l/oZqgSHZuQPBdgfDlVzqzSYPZI8fxT/4BT4nVXZhz
nPR1N0MtOyBMvoXiXIm543AvxE7CWRSVlZ6ykseLMXu8C2eXbYQLOwwqQFjmr4/rCrXaIFNQu1Xz
p0FaEp+it/Eg+hvJyyatN6OSYWjkmdNF82urEKl4QvydG5dREelRZJp2aQo7aqnNMsgT8I4yK+ou
lIZ8348j0fLuxvVtzSrB4tZinMJwyPWOTVdFSG9+RTGh3ncA8tfJ/ZvOvBlc6BYU8ZOde7VTZcS6
yXKR5+lARf+61sOCVGtq670MOPx2S6J+Lxtk7cXwtCoL/xWMbBnVDCrKRPAgSLyVNN62SlEh9t9V
C/AD9H+cvnOaJEpUPZsMXkqbLlnQiaD0mlfcKyLb36x41sx2ZzrABnrlpRU6Sfh8WGA4AaFG6Hed
BU7UClFjWxpBqTRn9Hlbh65Jq2/Atuq5g2I4DH1e5sliDdLBfhU7RgnunINc8g3m9YzvtAAqS67k
3D/4HIpbbf3oORLUAIFjVGobwhKsJphArqI5jeCi94iUR0JL31nXB9Yfjm3hnxJGTpp8p5zKV0ak
WfQxht09gZkbHGRD3Hb3aPBJ+uh6MFI2IzZwKL3ewCWSfm0QLgMwq+gLu+ofjhaNConDYzRpYF5J
+8qgDENy9w+NuJUEb1JIrvfWm26AT/+cdt7SYu9ol6/R8yEgBFPzJqGVgYpr6JXB0pyFtMztE4mJ
NV8K1LI6sKFcTDcfDhpG5PwfDg5tLaVC39T7FckntBGgAxfrg+E+Dwc3kPIBpVOK3DrBFJKNOnNd
GCMqHmTSqiZfWWVovQqtnZuaRZwsNxQ1TI5Ttd7XF4rK75SxXE+IcKrSmKZp/1YaqifOHgjp1zD+
rv71esBwteWfdwy42hGaxKa+xRRqwl89J823SP8GF6tyUsfkHVbaVy+gAp7ELbSlkLKu3g3kiJmq
rjW3LslhZU2Px5Ivwnpr1tKKzBBesi6FbzrKyH/r9YhmCBnVPE6gbG8vP8N+lGyC1UJ1AvIh8/VP
sC3L0NV+WsjkeyU+o8IwKtCOFp2t/F6Ysf6v4N/ZzpBe/84X5dniTNcYZHN53BHHrIlJd3Ni12HI
aiiNDG9+Bi4I6Bk/HPLQWzeS80fmxAEU/RMmf737YZGq9OUILvON+jjcANJRlFiQ9odC8UlN9XWB
ZDb8b+bhbark2Vv1Hb+yRWW7mpiZKyyWCltZndA+DWXZ2kDRxXCo6bDeL99BYUbWxuN/7oYfad3L
ywxVYhSvjf290VghtFBx2QD34Z5eUQSvuTRFKtmpIUoofgvzYocVMcgXr6Hz5aJgJfiFbb+q2Pdp
RWUiZuZI8B6EpK957ICPxObAtfcfF4zJbXmFBmiGHdItLYvpU30jNgzJurWas/dTys8ZzfsSriqn
6Uu1I+mxPvnpAeK90zHZNu2eAZazJUq3rFUSHJ+MDHy4Jxgyg80ORQjVr8uC8U3fPbca4HywlmlQ
9u25A4xeXVHEPndH/9YfyJnLaI8EqiRaTQMJIBB/IBJvfgjnm8TW7yPFGTPQjEBQgf6LRhio29Qi
PpBPcJkNdmtg2xyoOtKWUNt3to918Sg6crk2u5jRCIqVCZRvH6C+dawwSSVyMe+s/ZJ3/oPCaH4S
CDgTu84m52G+JeCIeRqV9arUAM/bVbD2jQVN0D9Sft8aTBdeauX50jNAsNk2tD4EZc2FuFrx46iQ
0/G6OFSZvBdCIHVsCSxteEgZ5U0LoKrArcN9flzTOuBdjieaN23mzY7L6F9g9b9qosWqs4yj2NTF
18UtfHbadThEHMc4rt1TydZLBYltWeR2Bu9kSuDFLG02N57sx3kDNvRmiBgmQu5PBSw3X5x0pjBg
71qrLHcoTufK1cdqnzHqfNZu5KGw8UO0Z82djUqO8bYcvnYmIRy+kRKYZAmgkdUriQNBHvReHKAL
3YlW4rC43ctlF1WDNRRIq4zAbVX33CGe31Dg57pVtsGDRnGrWuSdWbXdaWxBbQwYLkXPeusJh0CE
CqIr7LL8f2SQrIBo0gVU0Hnuyz2vqWv6kLcTyEU6rhGJQKbF+/nuHFB6BBe2pYGG7aqeb7eZi0Ec
50v0UF7E6vHAnMg2m4LPHRg2nBcB+4HyafwVQuu9ZRBTDCblKGQxfmRGMZbF3jRBGN/835YVeeWy
DiaFinaxt6YC5N2DBzpIcVEv93K/z7Ws812Es3Q/DIW0ly0ld88Vzhd3Y21Xn5HQinn9xkmgAi0r
F3uj8dOw05ghEk6KEX3RdJiEJzygZAQLqwBnhmdenSbMOAN+7TyOfZxdhnOOSGX40je1kBW++LBM
QL0kli9MZg5ZKPkAwWoCXBcwypCAKEYdutuogeqgE7BFnwrhkpR4J6+QC3zY2M+Zja0LM9Q1JWLq
b6ZH14AB/VdylycUj5G8KwSCCAvUbk3YhX5YeDyK8E0PXA6X4lUHoOO5J33fn4MATttzDUDTI0nI
MlTVX2yeCM1MblZOOjc2Sy1swR6JbhcPDLBXV7uh0YxzAwqNiXpKI5a8HXDFShnkc340xjjD1jJt
8ZX0Zhx8MgpaA6V8Je61bVCCA2+NoLVKQaxU2p/g1HXW+DKEyu4fHD6FRFevjjmEAIn+xbwIAIZm
beCdIIQeAzppzMMNiI5FrQ53bg1DvM332p+RuI6SWXAeLV7dL8NHbS7PZ/rTWmfYuwQk3/WN1KOD
QFiGaxLLJq3Y8IvBIpK1S4sWmGUmPNE9VxwnOUYYxPSMThbYVtjQiF/lppIVPXqnh8Cp7xBAHktL
SJ0n7an9XFRkWOA189dwLDAGioti9rnEIy1UcBxuKdIl/4jxglSGUhgBtYHmj7jymYLmXoKZ9I6t
YldYSc02819BKLvjVP+yzKhmoPnHMNQZ6J5NIIDNXN+EnE4Q+qI4LCPjHw2m/x25Ni1sWlGxaxQi
AlBX1bd8ufx8GYu9jcO3ccg2NTpgDwsUBljBQfIbfOLd5kQacQ6qlZJJm3kRWmXxuW4Kq00JsI2a
tDHaXD0nHWK4ltSTz0YoaejJ1O8yq/AVf0uFDq6I4vrNuZ6DGQ7e5COVBJrlcc/YD374PtG+YV57
jHD3rJJUYHCePpCFc+UuPYSqSURC8nBiA5OZYhdLFR1H+DERjEwtbjPNcLIEclhLA4iXBmd+OrAj
HNMIH4jegr/F3p40uUgxjG8T64kXALCsyajNdDchw+kJdUbrVlCMkjkeVvozI40/QGfq87IqOMVq
Y4h3jCKj60gNjdSxRO2n4fPYMr5GCCrqRG047ZCDhLKBw35H6O2DKDH/Pd6Eu2viGBSWJZzA45/l
mY6W/DRSCn/rs1LfXlYzYenbFfGOwcn4gmVOKkjknWRSJfX5UJGO+ZuSm2OCY1tVNbbwFtiXs7rb
MhnVNrTu38htGKNY8Txlr7i/jPeWejSNfg1oH7rHMTxn36G3odfi7Wx2TIvvDgp/VWKJfHMJw2cq
bLCygJvTf2ZOu8sP/GpBjNYoNhyJZaCvAVkDmPxbTHTaKRpve+WRb7oj/gKi4xKADFLkZWIKQDnh
mKoN2wKn2AOEqSgYeTpM9PTpRdsMEZ2PC2qkhRzjc3q5m12Y+z2xah3wgdJ33PLDhJydBkJkulyZ
Bd0Es6G7T4PusfnI3WlGjjZ0CfGVzXcwof7X0g39+dfu2a0BrIcCLAfsWgjs/Hg8roYZyXdQlDuq
X51mXwBtPCn2fjmEFH97Zt+F2C4pcPKY7T54Pt+p7fMlP6mDrtHl+9Di/6txo9AKgLoze9Mi06bL
CcNjfAW9V9DyGMsUgvs9/iC5J4sxywNOojYfZhm/0Kn0Q00eidubotTnkdA9hBBSOAO+Uqreaf/N
JUx0F/sz5ysHi6p4tHQx2vdFWONlU3VbUx9Qkrl5JpfhIacZlKDwl0SVDJzZZYP9Fn+YzUsRUiMI
zSREqA3ok1YJmQ4b3iHOgnmJEQooxwUkckpxQzDZZK4vvJKvqdrWyIqEQIgOnhgkGkZXHVhm/rIW
OhyHwoC+lN9zbmj5UJoSBdIXpbP+mXSGngNxgd9M9ZR1i0vEbJmHZoSbRgBVTY9dLJypR+YF+EWc
poMeOi/Bsj94Y6A7KjcJoDiz0Q9DLaeSkVusS1c0P1Ft9eKjyBiSkKk8HW9Q4+sLy+oj4abmJBUX
wDwpTcumqi08OcySGkgRAX8CXdr2hvGcvr2HkPv5duI8V6RPMorX/pWXDY0kRyePoFkXFXItHkEC
xQTQY0qjTNUaKeB+NrnnRQIdAzpTPdAHZWUBD6eTy6sHy+4/k5OCUJ+OAdw5Do3+LTPEiHjkCJYi
QJLsQcnyMbXdGBlKX1zV2RNoZArRN/vDDdnwSjUCyKrAns3D/AbeQ0PvXez2Iu9Sne28Pgm/bDNc
FZilreLExUwLgVtbKfts+E9uVHv6qYs9OTV2KGGTOa7CR6x8q9RASxBscVXZJDPSA1BHHMz6tYSM
uCQ/zUDLqZG4AeE5CH8pYLBG1Qi79VMBD8mo7LFy/Op1OA7L8iQgenu1kdHTOgwqC7qsvPr4Y8Vp
gVVXCFXnqgpf72d2gTSXPWBqVI7bmtLBplM0AoTQ1zBSP/iJQm3dbZEqu1RHoUxHqu8NtyuYztUM
DsKb45Gs7Rlkpn2hLL8NJln5UMTA+74oCl+Gc1srTbs4a0QCooKbyTdD6M1o6XRrrgncb3QHHDNA
zCkdYZoAHJK5i6RWWgqxFvPT1Yq02CVjeyfh5bW65j/P7MtVicQr6U/5nUDr0ALIpGuiyeddkfKI
Lzd0+WAqC9EztYxGJzpALq7c0mvo932DhApYKjhhB4IaUldl5EMPFWkPj3suypYHOH+hnsiJfoB4
BdKPGiBp759BEcgkyI8kaHChmuz+NZTMcVljBjuXaJx86lZt+in/w8OP6F2Wea4X0IeJGrVcK0Xm
wP1eoa6+5wwtlm4HnzFkjrrhAgG8HSUCtqSIHvkyP8fQIKPqlPMy0Ls8Y3iN0E/REnP5Twa0c5vG
ojRSw7OjjoLyVVg3df2xHQnUvczC1OqZA4hcW0GFp1oN+ACw4UEWssnkFs9IeT4cRsgMvmDJNl3v
LOZENE/E5zG+gW7kS4CpBRpaUp9HULBJv01JP9ngXaYsZ57JxAZ2cEGv5J6bzcM1Zq4R/kRc1zPR
elwft2e5zkTuG8VAx0gZeNKxhge4fWlZ6nmp3a+OHppyzRzIJyK8EylOTcO2XM8vIv4wDShfLGZJ
TPGE1LucVio4EAgK1nleEA/MaW5JLfv92KveWmbCGnNjklJE9L2+ornR8lI88em9rAezj8DEFHvr
wezKClE8NUMfyOr8DdAUFz8NsAmA61WqUSpHqDQEvrRZbi2g262uKMQ9t8UeWB5F7IVJjjCdEL6C
+U2/QPiooTSYu0UXqMoI/eFx/bfwFhWH09T5EkdWY5NP/ZDz0F/1eTRRXS8SfxiD8MU9LnUS+gja
GeZ/0bABiL/YY5JFDX9iT9/eRRPYvpHCL8MWcUW8Dw/LYvlj58iCGdevRD9OlvFQYGdGScxa1DWk
YzUFhPnuXgErQjVqnrfbjoBBz8gSFFCdejXS0jZlPbgJihekPf1yE1OPO+jAkOyE7GjjF4rUQq9l
1yxfodbhewXODiIlAKmi4BLffAAFpsmtt49bPETfoZLh7fvwR1dq++sEtu+1gOZdWa3tARQ3vssD
USgEtMP+UtD7FUVW6rhA9NXRKub6UtsA95Nx5qMlKcPgWOtwUhq7FhDDXMBK8lKNvsO5coJac/NK
cjYRdeocVwxgZPvM90XBEGc7vWkd9oWRUqssybVtRDh8agsA/BOJcXEyWdpoWCKomDT1W+ONhhGD
MR0iCTv6h9sPudmz+jvz4SjCdAldVZOoPOK2J+0KIY+B34Ka+UNHel8XvMGAhPyar1TDm/AdtXgw
kE6sYo+S2hYCPJPkfbHGR3Ov2+sWGNgZFLZPi+ffc69PfblkhImEwYFOyt9SjEkVbdgg4P9DB9JG
kRKGWu6KiX9cpqfIJMVT7vbRxgfnkAAXYTi75a6Cz/MZUnCmOaYwJpAOIdgxPfzjGn8lLIt8ArMZ
5kjSVga9QvnQgN01QVuwQ4rsNimQ2MN6jKNCFDZbS4K5iHc4C4oQoFUusQB/9Y/sQXbM8XiLyxm6
CDPfNSkfsGUUi94KapDChZ7YcAF8JdV3nIW2pvMZw7ifor4RT6lM8a8xxbZnTCQKl9Q5r6DXlk8V
vVcVneX1N5iQfpQjMQgmf9KRUS/xvS2c+TSDEpbuZU0HzzUu4yBcdAKLUxk6nEUmTADbbiJffPe1
HDdhPc+VnX3sI2jGF4aai7pPEzTl4ulgEfv+tAcp/Uari4HsfTUDzEUldm4EeZtv57n7TgyMkcr3
LQY578vkjpoFQvcdMaEI5wo8bxSZ6RT09x0gCQkBZEsOeBNd62EFlso5a3ckPZb8oeLBSfEPxrju
EtXMqR00XMhYXuFJojzp9eSbFieui6qloFa1z4gkpyVOZWQFOrJPlHuRKPEyAuOm1DW4/q4aRqPy
1tM9gX0sI7e/xr9Jb9dI6KF2s6EdgEam/BpLMEP7LuKknBR1eAb6qzB6pg7PS9o3cDqEijxNC6Qc
t6lEEfEp4FyffkMITqC0ZiwUe4WI780N5zJBLuETK/A5VKOqv8M2fHa0xag6IgBgZuBNeXVbKJDc
ymx3fYq6r0lQzN60jigMp5dTwIwAoB4X8v6Xk+u/ULMEOH/yPRBidIvGeH4rG0ysLj37MrhnaXlX
teVOsQtAtr7ify4+7uRDZ0i3VaBH/O4A9WDMGeQh+5zeAPZgMbEwJf6Etlr+3w+aHWSWwgOIJoZR
NBmmmEc0K3HfNadgSguWr6dsR5polQYSgXueraW4PYkW0Liia/g7U9UytbnF9NeN35cxbUG+t34O
nNJjnPSmZMhrnJKaZB7HIaEuozeVJ21yaVss08vPEnQh18eUeYLKvSD5QO7BDpT6OrjJDiDxFdV4
sqkHqUYgspmjh5rsXKOSdMrpu4l8BHxCl0lwa/KAkY2ee3xh+mWYk6QBGYfWgTzdNscUmcdIcnup
nKH9V31JymRrKUcdxapV8EDrYP1YRoCgoO8TNauYT/zw7RzXv+y5qeD6VMAi3vcVLpewsDPkmvyX
k/rq07uXYGo3ioomgfVYIWkL7H+EadBl7Ing4W7iSB2pwQMetMVZPJ3v0O2CUmbUtUIF0XOrEX7H
XXnoBNd4qOqa+ECTRs2hM9BqidlVHpBdLROulOFNmCPhg7JFSdqk0/IxoHqwSv/3nUPQyXr27WA1
FRPc007kx1YbaDqhL2K97otpLZ2c9ID5pOenlcEDAPZjuSAmiZ91MMnPRJ2GAd418PmVjvDm8WXj
oo8rEnuNuMy2p8SAx7iRt6zwvSLpzlZ3L5+Vh7KMx+uYwKdA61/MTtmZtyShAN/n0PKldFJwPfGC
6kyqTZCSfG6DskIzLhwea6238ugez1rQMZsiLgleWzwk2a2LkKcJl0Ik+YrPXR69rkIpVOIs5HXh
vhdPmqBTGKti1UN7j5Ga5ptu/w40YAu/cRYb0nMVKQfXnpvokETRG324kurkvkmrFK6A1JDHYMyo
hSu9EPMzUShkGgIU8U0ldIOAgFXvGsQ0B5/zQUJmc57l9RrRh0YBwUqPmghuAE0XgbZAdfZIMB8g
4BQUWiKSkQOWFqOjTPqTZFSc8U7yvvZ5G/RpB5yjyR0VR4zCmrZFa8sEGjJ+iTjaGqf7s53PCb5E
RoIZb2CdW1LE7HckoGN6AzMuazfwhWz6eFoXg1cve0XcEtkSRI+IdxarwxzJPRJR6MriSGGbLIzQ
ZnNJqe5S6tiDRlKMlGxpGg6hLTFCPbuyqfS9XEyXv8ZaVmFiHX5+v4rECdhcmy+tne2vcnsrr00P
nwBasZ2ODwBcIijplTmLWis/H3z7Fsi7uUvQXM7YhcxgkJqpjX5/4rd/a8AWPLUwa69OMIkH+b3Y
miwbLiV4Q3qBsGXYFbNC73M7kyZt3awZs1CWRWt94fba9be5fuKYojmPi0kF+4MKAnp1Lhm4VLf3
pK51EKPApziCIDXQI0MlQjSz8C/F5zrCGVaTveulq5SUpookAJ3F0V5p6xthZthF9KSm++70jF0z
Q5246EImjfx9JUn7lqDspOn1o27fi79W6MwkLpXNHqbAEpe/Ygx5S1rH4iMH8KVK8rjlc1dgxut3
udE9oy9VbKdn2MP59p0a9P2zpig2afe6qX+7WiZKUNPr2RTYDNSBHL2iGSjpivWrQX0vN1GJEzlS
zP0kLuIXC6juziR8FdiiaCTGVYOyMdGrb/6GIVArsPARobizyY9c18TFY4YJkiTeisA6jPol+vIi
3JaLqk1l+1EDRJ0GgWZAYFUm3eGYiyvKVMVIetqRz61wUvkruRsYaSglp7P5u+1sAGMzsekZ0QmW
K7k6Cw2z8h0DVSCHJ8OBjYm67wt8kRwZRnrtRuU21e8dgiIYFG6eiTCwE+heaf+Vp0rFx9y/+jpL
nMzskysFIURmQ4vcVsJCgTvyTodmrCvAE3oUi2h9jJPzz8Ml4goy0/FJVVJDqYPRyx/ectfp8VTk
WkmDo4lddZnfVU2hfr9pYhCDdTIgkV/lu07OFsg+bpEGDcwwT0vJUo/sWaJyA1wnw4cE9Jm3B5aG
TfKVO0tOUdPPFBRbisx3p3DNUyxyO90NDilFaWDiZ4LUinGKhz2s47zH6JHtDZmSnXlR2vHqYSbA
GKxFTc14La1j/Y611qaAgK5pmf4l/mtu8xbl6xBoRUjp/Dq2aNTIyeZN7W0T2/F/mywXQFQl8wyY
vh57PP7blq2AAf/aKXaYSWxrdYCGiNvXaQdRcERx7F6+ubVtQUw7LpZLrhNIM4kgU3QL1kr+fIfB
OsPJQrOgaxqENyYo7sToLc/MAReOH8BdLVkwpm87bqtoCZP9dPFt8MYle/P95ligQPlpLnNkZ4aJ
WwBfWq93TgqbUWB9ARmfhGp0UtbMKYw7e7B4d8zESlE/T3LomITFtdzur0JfSHn2IvF3fXgaLZK+
QQ/hTMYJmEqC3/IjORFfSMBooIwkiNnsIT89HvBroGw4I6zwK0O5QkfkyAwxvqiLTwsDM2W01KKd
Zx+20KWw6JWYg1gg4iN7QC0NdL9f6l5I2UgTpFXaagR0Nvwg7NyK1bfWkLfipNG+sqqNZOp+nfpF
rJf/fy9/5jFxLEr6bLQDgHV6+K61xdD+S7137iBUTuWqynIs0XPB1y5nA1RKUjVLXoIkHyrYzzVo
3R/3RtPgnZJ8pXo/QSOaB0vdPqxt86D4kC+RYUgPSwmC+G0EWh9xiiFbe3QTAyPwFVAxL35XsSLi
eDHiM0zRu6LmhyBclms/xL/KV/uiVjQwp4CeHMfsUkU0uzr/34+WLgYpw6RoMOgs1+j4XfxYCfm/
/qdw7Utf/6pgvuk0EChienHCBh3R7k5kSiASBCuAYcdxngjsD4FIMVtCf/yVV4ncs2JhJs5NKUi3
jUJ5lFQGNmFOs8o+baTk0H78K03xSICYjnFjZWbRT+B3/C7m7QI3tylVcNM9CqHMfnJdToAT6kMA
qrGwWtmBzwAbimIBDmRJeUjozTIrDddT0jNBpphPLUMSQxIGXXaFMtyl4FrubWXSP4l2uAfIKEDM
bEFtp+SDyLQ9MnFuyXaVC5r5J5ZKT1j7qQ/bFJMTDPcYkPLJCAVoqONiwrkuvaFbiIv7GHOOqKNJ
T/gfDiVGu0VhAz+zwACyFHq55xzTCCsNl0BiSkhF2UJihBFvokII94yRxzpPdgcOPx541jFzue/W
N5JfNc6ZrYZtelXzuUeY5FD++suvpB5nNZCQxiJpWsZbcy34d+EfyjFOOx29Ebh/Zz861VPOQ66D
i1xC/ERFgHybS6E9Zp+gmaKsvV3d+15HPwbct4REOvv8VTEuj9KAWrzJZSIR236DPTTsVG0lF6hv
dJrBPSZBdNu09+vmQ9foi+snp0qE0duoPyF5GL9nNWrySXQ7SagJwWP+lfi6jpcp2aj2wFPdTx5n
Phv3sd/99tpY2gmlXYuLG5EDlDZRdDjQhFEhjLWi8tXpxkVrWgE1knsvyLLNBvaLBzbwhb7Q/x40
rn3aegUOCmqBbFbTvnZBckGBNByPf5x+JSOrpRrfnUyBhqp3UzfI3k8EL9O5Am+exQ9iHk/3IyOZ
mIfqY+tdmJ4HZnUKdNbm0I/kxqWhqHcztAA2C3hmcQYf90WFkZCRWxDqYlEdSE8T6kqxvVjFvCfC
lIlCLgbkbrFj3nnsugeFFdUV+pQ4h2FLXAonq5m9nSCm2smFSMGLpPeRVIrx6vslRBKR6C4gDwj0
CH6KNL5EfFgwA8ovT/10EyIPRla6x116iqXkKDaxN9V/ay1vxtVLOJWf+GPRvm+1+F1nVQWjMEAp
LLYBUTcW4yEA22hB6ILgUPhStlX6bUQF7uOI/KJ+wWeZ0UA9xlUluohK1qbAjetdqphKPRvcNrHu
W1NWQbz2tSg5bnzFtcKqug+Ee+lM/G6Fp5cniBmcyoM7biPOWdHeyzwIDMtKzNaOLuorazNqoon1
P5XuWx6xTfFGLySvIrA1HEtmE+UcBwjy6QGACQ2gbvWIgYPsRCw5Oxu6ZIQ83Ps5ok6ihVmAqGws
eb1ZKDUIfCNQPjkmM6UjEEZAl4kGqbRWFQHluCPBaJMbLlT7MNMumEwqPtbp42j7sxJlpIo3ngF6
WcK+ycVlmFwZ8sjvSEo+5FIxg8lOOykWSKqAprs5x4HvtSUFf9dEb0zf3Yh03MOOmeiSWr88pjxN
/J1YHMQ36dBzpKwkRZFt1foX7/sLDb8ZpTSjswqyXak08Iq53dZVCDoyUvwkbC2LXtVXJsEhA88r
O4Yz72zCuOhBIQQqrG0XxqfHFITBb51RZV0U5IC4dTmO8Y/DdkyCIBBdUUEALe7kks8NmuLu1kFK
/qayLXOKOSQNTW+jB9UrR6+W5wfdjRZlNlYOF7xX4bb9SjBsqrHxGOskY8RCR0OTSegzK/7rtrCJ
fBZ1F56b8KQU08t+bAAJZr83LTYWw8B1yFqfczKTHoCyPT/2WMp+7spTcQPwaBMUjjrAMmghVjnm
DQMDGbEU9j7xVB2RdL+kw6XFLCYfq3uKhYG9YeVkBGfX0ahNWzXOUbQtJi7l0KUx6fkb3Nz4blVb
tuk0vSo+jglom4eM919Yg+ly2CwbwBQb2D27rOgXyWrVLoifPmHmWSCEIh3H3wIo2i+3e3SDQIwh
vpqnb6dSO+eQXuTsZsKTlA1gZfCPu/Gk46GiqqYByrjBPFoFnHmApYauJjCb+LGZat6EWuUMzqxi
htg73thE1cM+qlN2SGESMgS5Chtc9UbcbVNEzdwFggHqwMKbm6s7Qi4lLUoWaD4niX75tKtZFX1u
V7qx99o0Otwwq/Z79xEu5bzoqxSLrJT1aWM5PguX08CWTRi6YoJ+UG1/SKsqrITGCP7iw80pTRkX
u2ZEyU7+7YR9+30IQ/KmMqKZlVavqejnavl1okkGBcuTmWj0w8jrtf5f4/0twEIAZ4zuEJAzqyyV
f+xWKx/IqwB/E0uhuA80Zqx1kFMjLH32l2YtxKlfCcfGpaAKCzU6v+WTPjtbz2buLGFqSeJ/aKB9
lU9m8LC+7nmfJ14SyTb+tybQMcd3D3tjxxbatTaZ63ozkGqZwVrdUwPDq9Oa+Ds5gexTFBFfRqRo
ey6EZmKbS5dx1Hkirkwmh9YK9gU3JpejT/S6O6EB34ka3hCjpWM6IZ0P28VDfbwKGWIATkBiwFx5
nFoLOritIRz4XSJa2ccNRJ195N0WHLCjHU9OYr8aIIUUST/HnH5HAgwXYRDO/iCWyOtN4ow1glOJ
/PQjhjHtoFMEPjtdSG7kPZsqjI9tzU6zkTWqpRVgS87lVZo0ndDC5NxHAOU3Wg9oeHnkCRP/HRpq
LhuCgqjMpj7m0asRi0fTydIuPV3351G+kN7NujsjxMtQmM5bauCMwhzn5npEJcB58i9bboMOH/bu
06lx3v31jCSxR4DjrmXVdpywqVv62Ujwg21Zj1XQ4cjKyyz1yD3NWP8rr3X45NEpboMXdmx1rBBo
/YvalBgQBL7fu08yXvM3yFimLRXC9E97ayO3Ip4IsmqMXE9jJZiEhuysk1c6evXq1uMKk2QGFvIo
hpSX84ta+zM5gn1q3MpWAf7RaI9Z0Vr/aUwstaeqszIvUTqRRmkS1tpwI3ecfveWBrOMJ5r56qRm
xfzYMiqR9AT0f2Vd0F7iQjWUSde4v7M9awRgC9kHg+sFSrvG2gEmR145pAOvnesUeF1WAOoXfXd2
5XcQgRiWUFRJeH8njyiX9G39jtU+CdptB8Q2UA+rj/BVuocg/DHuLbYCKATJwhYlaO+sCO10hmjb
PaRMpPVyZHWbekvYelnHuLGpMyJeu9arzsuLbhqn3SLm/F91k6ujh0rWb6/Ck/uoKrZKmhaXek0a
g52kb8WJRVISBY8davaI9wBufl8Pvq3SYEd3PyimaW5mSc4WhzU9SRBoS6Lmnf7LRLj2++iFE9u8
DLlulkATbfJp6nXJ0SQdPTkv4APQP2fG0dFW3seaVkE+3ATDBNm9x1W2sgUFcMwsIE+tcFGy8MV0
qPM5nTpJm7cjJkNFYp13sgT+0U7Rmnd8tUD1RiU06JMmw3ijTecu519lItdh2bxVAe5Yjkt5kOs8
whkENhBgrCd3NG6cqb7nwAjNAaT8/qIybTtr+7QQ5i+p20mLOY2qYnn1oAl1zw1RwPDPfphKVouq
qvfm1D/BzCIOn0wXdfyi9DIwRFoKf/e9rogRhxpDrO432s7joeW+64FoN/QTacFDd2SmY0U2dEjn
ea2/+pPJ0TSDMPV/ICxuXVBdYpDQr9sBXeOeN8oSR5C+sLVtMMTWPWtHJi9TrELh+XECjVpZiRHN
A73ED7TPQiVeGN7ONcRJPVby0y79g1WAEEKZSpPy8EJRlA60Kynp76ZtoQ5KyV4cbM7AAFKjitwa
xbvYcMuq/GfuJu0f/ZzRitLzslR28Nrvgf/z3Ccv/0Z/4wQjrOib8AtNe2C70KY6SzPj1EHxSY3H
WA1Dtpad04klReimNsdSQZbRUqn+Qwb+Runwlule/ffzW+dfdG96NouHiOse/ZJoGZHRpcxhqdhn
FCIHl7SKRBEw1tXFLmBxI/vtZWNLpwnJ3P1nUWUD9w6zBvG0IrrlNrfxa14uHtWEfdE6rpIu2ilc
syDJsvBXWy/KY98HLhXAEZdcg/6KIcfz4BjXDlbvJqznHt/YJcNE6nLASXdcQhwawQvZgp3xQhO4
F0eLDIv0m9Q8QhyiCcAccD6ZTcLHgFY0ZPzluIb2KeHW8Hmg2M4UFUqlUB1A0hneqUDI8fNL690L
xLz49eDAZFJ4nrI+0BQuGnln1I27aHm/y0KA/rDETQEMs0nDJxa+mhfIAQcd0v8hkZVIl23bN+TD
bFifKvQm+ijTGhUQaw/eIaD0/fut8XGEk6VUdZuDefURh2l63j06OnEH4fvoB42kpb+h9OLbCXWO
UXw2Uss6EeruYO3vOfbwreNSrnStViUs2XgyRgeygrCvULorA5vYIzi0hvLSeH9QIFi1PtrufqBq
ZbT9qPv/Lf9oqOrpj+s94t3NiVGk1gQZ0UIfXGTzRudZOh74pwrXWpRyknQvDKi2gB4NCEwo8xCk
Btwlt1gocA1v+kA4GU6Ak7N03QnjyTjyutVX+yOgSOrhn/AGaiRk5lF7aiYP4w0ZKVezaDRLVp50
X5Zngdn+I71RSSoDzrc3DjZTzhjy/J+Zl6un1i6d1643ZImf9m4zQYiky6PKWey2F28uf7RutAK/
VmezmdtbuIKssFcycElGTVmqXmKn1B2vAdhdEvwVTL8czaeKqC294b7l99s7iOWrfC6bkqOQMUoM
6t25jeVHF2cyiYwZ7VAuawM8aKhnD8mvnjxdIsiq2C5Mq6/Mf0L7tPPvQUhX1mehonCXsXObfkFD
epLK9qOyTcxHUzd7mH3dPng8l4WNqdJgNR0kMToD29pCLXW92CIzAY7odAKSli7fg5B9oOBtt47+
JIWMFrcOZndUYAts8wg4s+2fCNs9BEvRp2SzeR3HM6o97/0beWJnULSHc7k3KPMijzjjfuRadkqa
Ahwp9WzQfEZvjzpnEtxMW0AxJMvRK9FQk/ZXtWiNiH01TceEUiwpIThADCfUtmi2fAUEfee/HsQL
/z9wTenK70fFa7DCrY4tEkGoEacfAzZeXEf+YwITqeIEh9dmBzoEqXC06cgKI0UnuwyCLHVMOsQt
QLV1FD9qGGwt89uq9MnC4wC+BSUQ3KSQ/hLUafhuvOuGzwC5oMq6M1vBy+U53uSNFxwBa6i/8SZq
bCbhSugjiVqL1IxbCSx4U2sw1o22YI3MOAcZYs1mZvzyGemjeIljCtxHznCqLSVyG7sBN8DBlPQx
rgnU+Hc48tuvVtlWex8tDjAhjszyrpAzdtlXEAi4xJ1IyeDvNMN60XhYEJOgtPX561sLGr9RWz85
WlAc4LWgQ5jxVfmOfEltHumLUHLkxaUjgEmD/FKu9f9zHYnol7NVJpGoHvi36CB6VnrX+3mh90n1
5nS2UrtICpXgANzjh4WdCihlwypvMs/XuuidkWVz5UcSajYn3ji17c8BYp1BqwEMqqrJv2lxaZv+
FuClUUJ8Q8kHMPY9ZrbIanZGKANY9YKUWEq8VAbEkfs7bC2d3OHb5+VSjv9eEDWf8Cv95GRkHy2p
GSGOd8vbRSQTDs+pAsL7wFBXNQYKwpKmPSMWXovgVFSTKZ1nC9Pf+Kh8Oukp7/rgXoL1QhHfPtYU
Gw3WwsGk6wMnkk9pm/k5ThOXiXAOWDh6+HCOTRpb2nBC56U315pBrlaRelGVup4sPXiDX3yR+jNO
TymfJB2bQUC1pwprEG54YJXOT7hC5m6AgZMWzlRBzrZNuPI53O17hnAbfO/4Til8Lko6G0Lg2WrT
gu7xUp6OL+2hrnFsJ/GMyA8O9mCnSXL0MtclV20vgP447cYmjZNv9AfiLnXQbJVC4Nim1AeDCcew
Gicpz3ZTi9Gsp1cIR8OTxvEeGjVEzbkd+6TJ0YlqpTM3V2fr4ZYuelgAk9UABXYaWydqYYKbFf7P
vfpP+hjQ+fZPpqqHi4oUa08DPPiStugkFeWPaTlIyo0ZoQHNkhwpMR6Q6eq1om+2HjrSPaYj5POz
HcAqbmwaSahk5rBO6tHMswS5I9TsCzjja6vUByyeoTXcCAx8M+YI7ujKG+mdiPXDCjkmVsIbYifG
GY7ktQmYm65CH2rRJteAv/YEX/pvp8Ktv3ruFzgTwl4uruf2hn2/dzS1dkCPJSH3yFhRnbobvIKU
+8e6oUkWvc9I57u2miga/nlQwdvptZiTugkQxno6eJIZXSUMNVi+7MhKtFoRGwG3R8SAuo3lVKtY
UNFDVVj64h4bSKE3cGuV7O94oU8FDsS2Ccja0EEG/F6wzAxLGrXN1o8U6VNQFIB/5wxxdgv3PAQE
T3UEB+rFPAw2a5eSUXMcyU2yaUwSi3UJKZqCguhNmX4QXO3SH+NrKC857sbmH2jJRHDylYhoXVN7
1N+kwB/0UbwkuNwwzyLfSSEf5t/sOTyQR3DFQINuIQDIov5Zj/LuSSqTXa1d8yRxMnY4W+H+hf6Z
5prqICxtLr1OEH4V+P+Gcr3xVJY6RemCXo6SvfuFqQTSKuviFj7YLt38EZMWpWHupk8V2eyATNyf
1ZQsVHmJSI1lAaG39quVCOc0HEHjG+Ug7pMxojSgjkkHNynXhfHaviB3+SFhOu7enj1tesRbkAFq
PWT2z6Mk9jtb3awYV6AtGVOepfv8Kl/tN8KUM//5zP6u5xxRD5fEqLwA5oMMoQBtOxvdxWie21BZ
kRn87KcIlUVl7wLgCWQ2/Aly++wRd0tRlSO8tKIQm2dfFRO+L7wpMujP/s9EU26f/oBHMhdzNHA7
/bhkJgb650fsaqhnWcwEGbXYp4XVwT4VOiY5qv9/FaOy0N8jHGh44KFQt9QsHTs6QDpo7vIR6jT7
yjYScSEm8lHxgbX/R+JhfdO47+qF+2f2qnOsxoErn8OmiL5oJpYXM7Qg+jXT7kIh5BXb9mN4bhMy
zIKgf91WgQRo/ysBPatVtkmCNCSuyLsF80bCoXzXCu2zaKhO/dGrvz/0IuMU6HMmCNxLTTLMHUMT
lB3ocMgiaO4hcjYVSnAeyEOmlZvss0NZLSBgnAszS5mQbAOUs83GrjhxBoV7Ul2IlCg2vczlN7SS
+65MiQxBjVuGCMfqQGaJn1+3Psde8jQzF3Cb34BBWYP0H3jj8BvBOwOHZsyJawpKbIIyj+Z5VD+J
87J+IroEYeSTSv0d5/JqVsTAmSAnEt+wNFFHnDw0KBELUgzoX8IO7tkQEg+Ypb98W6vmhmTz6FDj
iGLs2seBApcZOF/AX+voZ5S0xQL1rDiEVg2WfT9NcmrmKLJdR+rUTCdpyQYDnIHQEyoOJ3bqjleF
gvGNvD2aEDF0IVB59gABmiv+uGzYdJBf3xjGIBxKlRbDaLsXNJfZtZ2j1zVhtfnkPl4Z+GkRDuXe
His1YmzylY9/3F+CcOe6zE/fXPpLsrvjlo6C/ppi8PpwxaLIYOfUMmgfxA/5mUpVHoNly20rFxat
9Or/Pbf6jp4lEwUlfSOgQtOEBpYWEYu/6ljTDAglXybUMCKOUyH/ZfNczjViyLSpNSHV0r3f/tV5
xzqXyiQgUziad2iT01lFiSA26CQ2yVt5PjukATxZ2M3ll5UeRDwToMYMaLZbm5n974PU+zaZGqvp
Rgm403LuiaNe0OnRypao5Jd7sKvGss/4f88Byv5OhPWWGk9FY6A1AkcBXob3771pIH2bpCeqviMz
Xnv8eTEYAct9kISw2k3EToILj1GwfYaMu5K3KzU9ihdn3dKH/YZAOO6vVIHQeBi8CsDS6FUTuLug
2FebWEgjo/7EdVA7Jlac/2pP6Db7993SfovcdjUOlv0z0BK4W9MHMuGRnGcaH8/joEWzCb6k1Nbf
1kCarIzQOQHoKlCgivMoBvUC0Gqq3BNQnQbWebwMNcvy8GMi1yBuXuB6K9N3GdruL8cSkM7vbT8M
LT1uP+cpuHSNBg++hghcD7YFK2UiyObEzKnOK/n1YW7jM9u7EU2+4089vFPjfiJE5i9UkYlETbKF
fcHwFsrhXNr+V4q+V4xIBpoFM9tCVDlXYitTHWmJUvRRDdJbT2jELBmR07+BkKeXqvGdhiHrMlKQ
XoIMFrU1OqVOl1+h3PmVUv7OS5Zna/UP7TxuVcNgsStTKEV3d4L2GugyiEK0uWuOQpEQTfvEQpOR
qoTWP09Kef6/qrRStrN2sT8qCuCbXocteMdB6QscOBgwbeBShAMgntGRMeqWT46PiIKGcShfie+r
aU8jBWVr16eNC45rfXIzwS8aMT/GrgY/Z4welffzTuDpksujaw8VMHeF6/A6C0s9OGKCFHpqEhFs
C4bFU/OwG1uYZAdSRxUCZt3sbUH3Ffa48cARcUVJnTQrmZGnNd6sbIaut3QL9oJP1sVWEM4pHn4i
tug9d1tUfvH6xA/9xFvhFr46fDy5Q0K4ly4unoSPhtF6nQ8fvxuLOdmwabbC9wcI81JfvDduuCy0
jDYGXntg/Ve6tuImKoxniNkEheJrU+juDGbuI2XRc5lv4HEb6t8DdEDw15NqFtwpwOpWrrctInBv
nPYw2FPdr0uFbaTwmrBNc9ntlXRBhrhXWWk66lXg080nt2z4aNR7GVCRxh7OFyyi/6/6Xe2Rjmu6
hY6BTO7Rilx4ERuBksQQNanK+8lmjDgRd8lqjwhqMSsdYweEfXn8tqPNWl19s7EGbUtzNHbhOmYf
DYvPlc92X4YLoHe0ssklQp9aygwlEcXGbgELE5vKvNHs63eMQPk5u/MbdVz2JvjhbHA6qwXykN33
RZjR+VB7I5gqBuFRwOwctFN1S4Nmd/H8CYcAw+ryNH3p4W0zVtCV2RxcwuLVDTNCD9O6D5rh/5IH
u5MquBUxoFXy0JPbiWT2RzIY+Ep4nSI/eWfLOTCE+KjWSLxK4VHBX9BWaGso134vucNAokV5+37p
CxfwCl6jhbaVMkH6deBbjlYyx8AV4kb6Ue38faSV0Od5RCaiFYIVs43LvtcaLx8Qyn+jp5cZ3RGw
V7Wu9456IZXb+zcluksgoLA1JZzle8VVHVMXllRzz/H3GmFP0glMYZsCUP4uJ1Vh0ttK32Sjr8zA
HC1GyTNYNAyu5zIn/YZxcnnDhCxC18wjcOdVPPt82jE7wSqav6pHX+1ZZNTIYdsE7r4zK888PQ9C
y/Uwq7Gw1OvQLs6xfBXN/da4k+WQVhd8JiqAUzPx4A02GkyoDXVhUU/SV37M6qPEjoZzFk/yldYS
l7wE7XOlWF1cbvd9QhFPuGpMkYHh6XLYRU4qr6PQadvttcLjqlrhPEbzLKcO5ObAVdKJCjX/GxWq
cIjxAUNqKBBw1aviONM/jg4eeStetSSNNj3BRkZ0WprmN35I3EQ3++Mc5YLR1x9wu71O4AaCFdPr
VB7ZdH5EyBFX0VPZt6n4igiKFttpS79wmMYmSiqwIoxz4Bz12Mt4Cf4mEshVVIU2pUAXfv6GaV1n
zlcIy8/UjHahUHbEK0/ExZn/7Xz6cM5KvnOSOddpMZB85oDfE8NVZQkuY0QMCVJKEKKtQ9IPitlz
6n5t70ewKXxCkxMKDLlFLiYOzi3CuC/MnzXrIunqSBdfMR4FM0Hf4PUx6ye9PbcROAsn9aqnicxn
tnw81cyd7VSLsAII/6ut1JUfd2aVjMu3oGQJ7UIxG0Y7AYAFL3Fqi6N53APVaESfV7rJQFOSznzA
Oj7/WoGjCrCttdbvVmWBRXzWSiA/UtazL0/xz0yqiAEe2R0hj01BuFjVZqP2oSfZYt/GKuBHUVrI
I4qLNdId2VbzkeQroXK2erDHR9GeoyfDkSipkdgS+7LPkQRl6dmE2jVuFTnyVcVkDOQcmN/3vGsx
V+2vP7tPUgUwRU9Un6WrkhUkH01cR7adiZqbNpPLUsKLFhdNDj3CmQkS213zAEbxEUgipI0knj/8
dqjuO6DI3IG4LDWUljTa/8hh5YtL2Jv6Bc2UcasNeHoxMQa6qIvrQgVXS7Z9ya3WMfkHhJYOWBQy
j5eTkIkP2JIDxONS3YfyxjYP1rinXtqOUJQhz9zulxtUlHup6lolNyAGPs29IQIbSybPMr+Wxfxh
BaBRgo4UTjSm1TNzu/toRMIuwtZhGFI65UMFzYUhq7yvB4tD6l36VIcT1gQVrD1/qq/tkSESvnwW
/d7fkWrOTAIyqEUy/WV3FBeuAcrlubWSzAD5u+YZ17BdCfxwDG9Nf7t1EpKFV5xxzkKxhWJkSd0w
VKsoQSYhN7NxDdvqp2H92WUjqdig3YUirHckrCm9HMB6z8hcQTGFmjQD38XNHeGzxxXR3GrGd0o6
ExWpwx+AwsvXVrgfJTyWVJI8V3t485JAKpT2gPYFBS2lKFFNnNXMZI6CR0pYT36ZqqfBwHxnM5Gw
AxyBKGqazXdItT0ejslQJDt+csYY/DunrSuifq81uhggrsa2bpQ18gasoh6CK8+fjcCf3XAuL3C+
P2VIipn12hfHl371Edf5vw+UgoWX9q0Ny7NL7xyn1mnQrXi0nofOgINv9iN2MSWbtcGRZe1T+8WS
SvHn78u/oFnPo3CuH38QuGNUvVmI984ez9HTZ2o4NRkS19BMWnw2wTwnIQEzFLaMsn23cFOcF0u5
kcNMjJq0slapGDxGtWC1fV9bw98a5mGbQQBK80lm4lztyWonkptYZv1XvGtZt1opxp4Ao5BTFLwH
uTC8aKm8fS7xhPcwnopPY/hHW7dsYtHd2OPxjvZEW3tZ0gIKYUlaVZp+K4hfrQ3WpCviZfSuZ9LG
Pi7ei/+d2NKZoj0uv6ORPNn/yEQKokEP6SLEVHVSNNSl5KefyirDaGp21dJ9oe62q52JUNIGPVNI
6qSpTAjM9iZXep9iUpkbpNfL+kCJNMHW5s4TFsDY7+uVcNSPueCNwx90PSudIc5UucadZU8bo5nF
QbiZs17u614UXW05zi1KI8ogYy+rn/9940ZrHkcNHrlZiPGyUruMJ/IMNBpdPUJ7p1biawvaMVS9
WLaXD3eKykEX3ognowRHbAGVyoHhfc8HFcQ+pGzMUEmDXGNZ3jOeG+lVlqAH+NribzOX2cYjcUxT
LbvJ5qpqNQQrEjpjb1a4iMIDkNYaKCJCf8JcA1wn0OL++TWSok5OBmTgGUlpCOFsqyw2bJMonBxQ
C48BUECgRzluKMkEavyzgS6ncflWVXzQT8EKzlWPgprf5pPVn04VvQ7+AgNogiL+k/rz9oZb3+iL
d4oXLptVd7q6zezxjvZK+YnAzGSAkLM2ak+H2YJQ4N11QBYLkXgkEn1s+fN/k3LR6nsMkwxcpzbe
KtWUFHvEAFwic+6Ci0sYqXv2r4kuy2z47Ag46v23YFverBIxp0UvPYvaKIX91mzYCQjxMZ993I3P
ooghmJFbw6HWmoEQ9Sfcas7yk2HslimGS6GtRNqwrCGGjMJ8SR9IRq7/oI+WAKyo3Zo2yj+hyKx9
Q1pQ/xaxylTQn3dF+1f0/lGTh4lSzYzoN59zM5oAeLxlHb3huTcbwmO4X1v8sqAwzgrLDSGSHN5y
jqZ0TkcEjQqh6kWzlcWlwCAT1FsyvdJjSUqIHy+T6ucYlygO2ASZW8wUOgKOMKp+uRj0CGQlPpzr
N8jo9gu41fzwxvo8Iv9s8aWg8mz4kODEsMtspH6lyPQ15EwTZhuBo1WATouXhWmz8X3pV7dxfbVx
i8MWUu59KDHCebqatO0a8DfLw2b7mEO9ekPSIOFCEmMxJgX589qjWrBNAsFX4KREcauWJSEHq20C
9rWllub14hnYEReiteg+1gyKLuJAnXxRX4rl9IhlCZ7GRkmX0A+/v7VGAiWD2WaU26bOsTwB69Mz
xNtNQsj0BFxR27u5Jz3QJMC1Fi6ZwNsONvKjP6JbbeYIpRdg87d+va1Q2MptVB8P3WRGDRZirivY
mUOoHmSH4J/8KqmIMMkzgZCYf0aCAyVmi7BCvq53DyuN8HiWcA8S5VYfH6I+dGfKn+7WwKiyH8B3
KuPFAMUqiGxjMRsTGST0YQO4AWp3Qkd+HyNW/NA+rl8l8HFjZHdHkBHKJV9bAisvXYiNK6QYuTvs
ZHBFo1gO4iWLhLFWi5grtmteHJhesw4xqk7qbix9KBY9yQYDiwxHmOocvXHH7EnVkGHkusBJ7GOz
SP478OwENPtNEUz/p8EZvCWHxk2F+n/nnS4hLYo6ynFEQH2W/8xXD2RicwEPmCTGfOdJn9lW+GIl
fcf5QOuTq9nTkrYEQqa87uOZ4v4BXuRIaA/dPc8OwKTED92piMx9lrjjWfyCh3y7Im3Xa8fTpmhu
bRg/ECMdqhseQqO7pSOvsZNnq56mEGdvecrPeFuduvrXzz73j0a5cUS5iqSCVeJTH0IibV4uU9sP
JBPqnzaRpNiGUdJnhpd2O62F6+XwUIzXYwNG47fMgVr7xtMVVgw7Ha3zfn2HNJM8dv6bANkDR2tR
amkXVWWfwLQy9kqsSNzqnkNjbxv0gTNTjjLmkvolVUqrRBcSqlymzAT57uDMksjNIIVyeqQ6pQsq
eX30qxWrG25O42yczqyzPtTpBOA6Z/Jop6FMeejOpmFoct9i/5KCdqQI0mo8dqTG1beLSQOI5tVI
mTOGasVhOVdigY0SFeC+x3PhA4OYFWuhNlWmhb9vBbgEQh3kLIuMPSeRTHAUOGtPgfCyfj/8Pjp7
3fCmEP0FbMLwMBcp/Ae0xMZ9MdCeHJUYUDrHVB34fEVN07cg5EeMrx145INLVSgGUETVRndvJSmq
Wpd1YMxTVoBJa/F5Duj6OY4Nb0yi9LMOFnP2lIZ8LkGIOCsFMVG6tA3QpDQl49S/NlogNnSWj5gR
cuvyaBWk/9M17qt2mOfGzt1zKqqNLnm/y1ckNPVrY3Ew20tjD9O6vKoSG7dDB2pvK3u3k392HqSR
bThDkouILfD7tRwGQ+85KHclKNZM8Dv1pY0Ew5YRXVHcKLbm1LO1elhgyUBMh9HdV0kq/lKUZDyP
xJs9FERtF0LgGsm1dhE/Z2prF1z/k+VE9XZYh3SkJpWvL1mzspJcSmrbQpUeMyH83lyXmFOUw6KN
kh6fzf1nI+v1YxlMZniDFhL+ImVVsSx6eKGK7VU7UUkkKKK0UKvB8bdzdCwHc0IFR6nwbwH5ijcV
rCBL1Oaj6nxrZLhkaeO0c8v6oAKoQXXu3axdYhaCcHnQRPP9TWGpxJJj2471aIu2RRQqPhSjml1I
a0c2Xz15X2Duv33sY2krPO2NCk797/XEmkATf4R+ILyi0HHy6dna0/NRBj/e+vRP4FBRfLgNiXd2
D5cmdEJ9qBgMCLic4BipQ/ccVB5zCTQtnplonSFDO8q3vwfWcCV5Rg3wcEgG6jE88cHY26Ot4EXQ
AmmEmfbbQ5GXAzNX0cNEQGK3ilqfqnfNvpR3pQWPDhWAgfoJ/XRn2wzJk/lCpbzQps6yjcPlQtYm
97DGedsKueHY8Q6Y0WIV4yvBSX9W2rmdv3uHDNS3HSb3QmzmlHs2/SO5rMyjzcAilMuq3D7tjb5G
UZbISzViCdJpMPs/+f+4allw2jju8IWgXnKEjKYO2HtCmUV6Ktxjjnedq85ifJ5G5IuE/hnWDQRv
rv21LWI1jmrFy1wIklI4iO+XY4xYNUMjpogLQkIbNYfh1uCBsTxRpSEPFHQIiFT2M91UQ8J34lac
WOiQurheRtrMqk1AFdHu5lu41MNGdekkS772f2IXRvHlMjgLo5Hzub5P6q4LW/tIa6mz+dT1ZwLJ
XN10E51zTXaBxitJ92OQQjN3ya6ml7KkO+jGq48akUEsaiuDd0Cl3m2GHVcircKZzigae5RFVUrt
ZTlHxqzIdSBDNhv56zgXG6voTmElVchrmrFn/PAO9GLeKtvuQiRcdlPh8Y/8z9Mj51/QlWLwPVIs
IsJsGdqquzVyTbYDSMrdi3QV2XIq36VDfOExpQmq0KgNgIEjmw5PeasxOuM+T95ZydUU4ABkuK8G
46ohUfZfY+u1fkl8x1hBxgiDjLvyE9ZBMdiXeHuJU+M0UXkw90h2AcrRIRuTHpR55TAJj5MQjSa6
wJk8Vp3PzWlFxEPiPQyyN1rTvr2gEMGzVw/vOswdiqQRUQfHhCqBuiXKQY5MjKhfyF32T6JMr3MM
jfzuVtw0WgVBfWkCbBxl1GlmELNY3hRBHg3EK+rLoH/wDKveLZLtOewDYw1WiLwIniaWYLZB3RhC
7GUnfOwdZ9x6Z1MR/VfYZ0Qf1d4rANM+h4rtEaKmGiqLtdT7v28Cixmucjv9zTtFGxqGBN1KKvxI
Xr3N2+ekF3S0pZ4ruI8M7tvOW0rCTBXHJsMEyCcCOfwhV2fMKa2bgXCsQGQtjx/8LBGQFaiCdmZj
XA2XzESCKiLVX+UQ1z0nu10iIk0s+HQsHE+khDH0fL+jv/AMn0hqkLdLUCruUg1PoCnl5ZjKdefx
il3kvig+U8fj3KCGDUCju62Vgcqccn34h6DRXRlSlTvpg99eVNGjJIBeCFsWEPP0qcrkRmRNjiic
Yql7b9KamKdMojIJLt6UXfwaplq/DPeiLmU0/WrsOtwW+HK2n+dos6IDTj7qNXlQTrisiNrlRtg/
bOSJYdTZflm84lw8vzRWktWO+yTRpfNxCs/zQMvVUYuSp3vlqxpp3MmS2CA9g4ikXx0LxRtNitzB
u6nQWdwZoaHvHdBa0MYDgS3reEosexcUmQnZpG/ZEyi9rVj0h6q0C6QeT1eTdLptixxT3sY0twO3
bUUuc0dKn3zwbpQZ52tV4/CzEcCC3qGpWTD8ewl5xeCDvz/dTBuI6YBNITedyXr6xjkDnj0D8kiB
uUPXuwX6PjP7Ymh9ckWZa3YIfRD+y3GEx8/tIUVmMCxjDqNuTyYtq07PWekSTN7fuwNlgz6l6TuO
Vaw1a6Jk8EvuEwlrLevkKi6yUKhhnxYwzDjXsQF0XAcG7MS6+kZfaYdoiFPrF4RY3yWgnEJ51MPL
kIT4O5TJNAbDDWIhhQcV3dN46PDQ/VimpPGcCe42sp4vZml36Gq3afcTFYsxVVcdRip3ACAQCek8
ahwW43o5NQ9+vAFEWEqFAEZySm2qMiuBCptMUn/X9TRRe4TLQxTuv1qbwfRfVKX85MRb+tHiV0lB
iOW/r+uybrNs0xLXRemakV449L7YxYgt3NjFuA9Ut5thvlFe9Vovv1akBpY3ngG2ExDZ1D3u0Exy
VDjJt5Pu5IIthGX9Uww5hp2Q+0LuP01o45zJCbnIUHLC/y5f3E45CdVgBSwLIz412gTB2YXzlWmk
OXzeHgi4Yukv9qpYvqUe6bjmr0t9RI0rd5/bFqxOrhw3v0rmuD4Erju3RkUmEBKHqEq4TX1JmZqN
JZjy7pNsI8GcOQsSf+rleILlJ+FzHZTs5ZHJSIppUWRv2MgxpJEvXLFTCzASyr/1mD6VKYdZ5C5n
6MH79Mvc0gcvm6ALQ+GmVqBr4tHZgL0dXipdC0pei9ehupYm8upp+8/frzw1Xu5Ai5ROpxGI8L2h
jxWe26H0DEBar2utmWO1CYiwz12If770H5jXRxQhzWyOU9R61jRqwgrPwbfq1mnfqS8KBIcAxquW
YylSC1nqassi7/6kDYs4/AbnLFdclCI0KeovLJcZneEjN72WGiLpBLl8rrJc+/p/B8b1/9hsovB3
T4gZPPVoL4AXNH3Hbqp0+o3JRt7fPWNEV1xGjs1SUJLSsHAvtSJg8i6zgFwl4Rn1+HXJklKCjlYD
UcXueW6NVRZ5Y+POYOYCZll4rPGyUalY92AILFcpg99DFRpT+SmnyFexKCPCoOlmvSFMtCEcFZU8
3bOVOSmvXIeQlUZiZ8C/wuR/5yaboCwWZGFWaFro8Qfij6vYlE7nS0qGY1/EjWNwEEkzrE7IojFx
hslkFyeNT4RFnGn+uoyFbgON1cwR8X2mRVW8IWrQcC1k9wRJsSeLA2IeaTEube7eTff/6J9frrWR
/eMYdoK4KIaOFuUI/bAUGD8gcG0r5cR2ZsBiBG7oSrHz+TA7LT2VkTamHUY6h+VUdPyOl6WgqyBi
CLb0OIvgwqbXj7G2gdv/lKBdyFouc+KLeGKZEzdyZGAoyKVlgZA5lWTOnQik3ym3CI9h4caz7IUt
uLaC/eSC8esUekg+cp5mwcs/yTGo6qwkDo1hAroNNVJevBEGuozVzBcvU7JMTJuIIbDcvm6jfDwa
VzYkg/VbmO+QVCnkdmhCGp7LASR0Ggipx/5QlczUn1zTd6qVAsmzat4x0pMT2/s8SJT1ARl50m/o
9asFkoEojqGo6Yzgsdmoq7ay0t72iYVWXG2co6k82IE62vSkEbOwSTKRgiJh3lZ43TKRqI/lUMlW
moNdPdLoUsMC6nXqHzqVWUXMQ9lS/FFcjScoqZ6Jl9iTgY+OXsnDUl+jm0DhJAdESgR9XDYLjRlk
2fAQxeHQ6/lL+Pv036RmnHDkety3Tsh8NKdA7aGDd4EMv7oHeugl2j062c8brz2IS/Mnzleu7SIY
r5MMBnU/KIp0cxfjbaK9m14SfdyRGv4uO8dDWyIMFhwmmM4ZZ0tYNZqX37LbRlAY0pA/CCpQsuxm
oD5oEabWpMZXicRel6nzH45zBPTaT4LvR8sdxo5o+maK1bO1gbgtGjbmnCqGt6WzYqT8ul8N81Zf
qZkVxIl88j/l83yyKF73GjWGhg2IIm5APthRLCcbNrYy+bmDs3eWBW3L/mS4aAi1nPwMbwFAw6+P
n3OQJvS3duL8X0cxF+f4HIw/ZAQwhVlEUkBggD5uT8Q7w0gQVk642VDZsLBcGy7nHly9wUH3+dNn
W2LmLRZQPH6Kc9WULr0nZI9PTVhyIH+e0egq7ZzqOqUJ3fv9SqjgtSLgqFSdRu6b+7FQlVEEdWdJ
3kQJ+gvTjM5kwR9smAWwKTjx1OpSoJQabwcvgkQ95zUbom21zHXktRpLU+N3XjXXdaVEU2cvx90p
m82vssVsEzbzmIvhOtUNF9GG9W/MS7aEuZW2o5dhs4fhBmQWBAPY5hf3guiTslvwk9ucAjzA7YZ9
cLTCU6wVLHD7W194t8iE+Yi3FEhxAIN1SVlLyA9QsE0Gbvf00kDNL/AaFpPvmI7dScMWxUQnciT9
3sKFQ9nkRgi4ZQGSMbmc0zCiwSaBk5oVpIFbz6nutfHXelWLdIPukPPe17eEzQXLnqhMS9Xgxr38
qpp5f2d+ufGbNywUXKTeA6isXoCCna81d6ydXCnyVhLGuPpiMkOBb8tJI1vB+3MjiThpPUxyg0FF
XFKF+tavnckrpTRziglzS7D3qoB196AIfPNXoiq9OuK258NneN6qBNs8/YFvZ25reNXVZSVkZVNK
m5I7XJewr9o1l6tJBxlvJerEOExrqTYzvWfa/5OtvfCjw5RbUhQd4Lb5ZPmwiOWyYxHRfpa/dsmr
kIaid4QOEAyVNFd+mVNdJ/2UVpImEV0fw7KiDU6tScWIPf3Y9g+TL6BMgKWfqVb1p6bxEC3dA5p3
QUlNsWskbnZeH/hHUYZpT8aJ1orIwIiXlpLUp6iW8hRjpleYqCZtLTam0yIhWqlzx4l+Nu9PUD6A
Yc4catoUfm0JzR149qI3NVWyE7x3P5MYjyXUJUoXdpQXUyDNXihVsgnCTiyDCtFzEMSMVedB7Oqm
WQzYT1Tn/VUks3HE62VUIDA3fa5cnoWXXBUz9OqFC2A03jOWA+epmvWlzMb8jTASgQeDt3An2cJ4
cnI8agTJ8AiglXEsEtgX1VDx5Kp4w7veCcf4myVF9vNredBIQXx0qbDYAJiMmUu3YKwzitPk9rmE
i4iHqN4gw2INI+KwlL/Rvc43erFCYTvsA8zjse4ErVJ3EH/Z6aLkUnSJmka9WaEGRH9UsHzm/X6Y
tb3+B7Jlrzp2LoEBHhSFKJJV0GgrBKb0yciqkOYuAUx+d/iL8BQoP1rG+T4Kxem7jhuDb9lbmHC0
5erhqVTsfUszlqLcCZ+OJ2e8tI9Ds45ks6Y6BKY5JsSB1J8FTCX/jPV9hxPiOia+34nGNx59+diq
SKhwisD7DTRc2e/GUnMQCX3E/gUyILxRnlbCV0yOWno/vurFRzF8W0H9WN2zh12mlC/AT0TTGpoR
cNSn0vYxfSTciHoQVV32xjLesC7J/U3O5mRmiTC3GKgLdugfhbwlLoGXUG9boxE5q0qxbHyxX+lV
MLN/gJ3SZjQ4s4DtuEDc2wvBZLRD7eQ3jGRldLP6nRm7Eq/1QRo2BB+CE0KK+8uC0u9rHvPHBZ1Y
HyE/vcZZqhW3ntwQ1wH1MZ0T/Ll7XaHTt/lnXnDam2uReLeJHmwdJjg0yCPhpKIRT3x9UzAAL+YW
5g3GNgJcQ/re6dKz5PI6ABwpAyazmjTMMJ7lIPeusOnbyOSx597vsbafXXFBWIr7zu7RoAyhRVxe
KhZiRAlD9jinNyWZSnUJZq1S8XiGrGSTsmaccWCXTax7mOsE0oZ6VF4bLZdQluhGg6idXJf02prw
ELLn/lPY94s/gOHWWyUJAg4WsL06CvkJV8jjfKFpyRtTnTvfy7nO3eehybMnSh2AAH6rUrFxtuH5
XvZ7fg43FZLKImLAbkfcKIig9/O9ydtz6h18FYTiY/+bi0vYe/fML/9r1/JFJ3HL11NpZUBfvm1K
g1Um3YXL+jrReFj754N5fBvOE0h9wEjxjEN9Sxo0u0Af28nFDZ9uHuxq93nfO2bB4OWlgSoB4A/6
CvlKanQhcPvXwfhTCGP63aS7xK4D1Pxc+1vqeR2vq1pbAzMDcV5CggsRXw2Tk198i9spgMS50IcC
sOftcovgFqEIzJmzlxbV08N89j4XvI6oEG3/VJgiFL3rJWpM+Qwt59gHex+1Tyu/x4ZBFOcLobR/
bibR7OPfH9sROK+g3jN17XeJJgbLxC5dRXd15w6ZmU1LGvxQ2dyXh/gr+ze2gU+hQtVXXaswPmke
XcHaOO4rFVy3aXu6+KbZ+lXbVUGprgTDmoPLE9vm9H8ocAQFxf61vb53xN75sJz+F2WIFqNiBOjQ
zYmk2+yyfykuCbEXT+p+ThBAanYaDkxRu9ZHvF8tTQ9B8Cx720WhaA6Kr7mrZILCsVGxn5x7Asqq
9zG98a8iNRdZVulY6cfFK8zAL7Wm7sPYYajK0Iy9TTajrxzr10Ks+SH9w35K5ePzntPVCmq/X2kP
xYNTqv20D3zUj8VhCb+0fcYoR8EC5+8MY1TfhxcFk4S5HevDGLkBxME7amZA3sjavHq1DbK0d2b4
+u294bNdoZlEVBKZiNCVnm3PkjHQxguT/hNggqZ+XPVecqWk34r9KR3bGhaqoaGCe3UfJ3jjLwmx
iT/R033SH9YJcgnEI9EoMvVzdRH88NCD5ULRLh6VjtacghlGKLXDgLVqr2tMwlGEyB0imJX4V/St
/UZtVH1UapjgEh2DtXDAVISAfX+IA5jEh3Gvk/LcFpAhiZjTsZA72ZcCWEs/Id2LP/mfLUyVPo6s
27D+/q/3qJStAa0uyM6rl9bAOwjzOehiJy2UTNWpGRnMuiD0XcefpEs+LVhdu3uPOOdEnJcmgXMY
q1iUYUTgpppQ/zvMH9xaDTRHUpbxM7qwgNl7UoVPj4BErKiF9B2wunIqJgW5MT559oq6knu4s4Lr
BD0iVmsSwOyfCNKEyHes4Qm7QnQUBTCb+/l8fn1tKgIZlg5uGUoIsdGn5jjKuk0/2NDpxnnWAfWf
y9dg37dASEAXvYefh0WPYkrx2q/vGd8Ln6ayrEGzoKFni5WOy5LjoaedPyuzFJUuFrrld9Ymzo7s
KIYa87VrcEBFXF/U1z1kE/XLBmly8WK6mnIY7akCRtBB5KscMNw3RT3WOB5Roh2hilo1D7AqRUpv
HLgK2AJHlhz4j0u7c1jdeim96sdWGVIHIqlyGB8jAAi9wh2TNsYAf04VKSnlpYbwjxNVQt2l0Hpr
XCNkf/Ckda/dZMOmHWXQTdVn3KKjPtL/V4JZtLThrVfzsmyKqHzFYPfP34IdWiUWHpsDLRkXpem7
Cf2u92djrerHgllKJ/AYJz3HTTgJHnXyaCUEso8dwNHrfcPez7XJyoefVEwnsrTPn1HDvx8YtBTU
qJXe9LyAzlSo3OhEcJH3hnhJJqzHp61ZPwH2fVY0jvdHLIpGKhs0XyiwJ90qoY3KDzdPKM8TTo56
f/AYkCIslj7taUlRbLbe+xasbDWbzy1xCoOdw8AgM0ihAwIHx1GVJgPQMN2GMQKBtSwuyIod9LGH
tFGLYC+AxI1mOrB4hh9PlWfA/+cZbDAiitJ5llObq/cCgW02e2ZZ8LsBwMra983I2IV0PpargsCf
GEU31dEZw387a1BtYOIFoxIkojhhmB15w3rRmqw+lc53tJeJKSAjRbuXplyEljA4DKgQdsBEczTc
gHvMNB4CAA2pBtPZghiFLHfC5fh+G4RmDYV6jGeq7fFk9WRs1iwfm6dSqKinPP0SZty/EsBgFhc+
JfQ8q+xGZldCXhdRuN+JY/iHrUjyeft+YLy4krI5TrD1bC5wOSUc+Ip2CGRl91qyF6l3TvRDvAzp
auWA6jOyb/9km+x0PoFCr/38295UUCNPonYSNvz0x1rQYflwMCqcsAVLiWvTC4Xv5AJmYVAawfkC
whbReujzapFcN0rovBvNFh/bPe+DEvsHKWIDpBnsxDWcAoTymGvpA3AGVgtY0cnd3AZte6xea0c8
2NiKYMdH2Qu6n46tIjCOs0dNkJ3nZKF/mKlN0HxmKOZTn5QdcDR373wLRrb22zrXMYanptraH6VI
69ehNfb1ODJoMhYqIjKy6OWDNOWmUlOcKXD0zYNDHxY/IvqpF5Wjsxup30JwmnaaqQgd5TxXqG3l
59Pm7At8tWa9gn2EXoz+DbiPto3lGB48WokCgtczXtoXX6IP2EVJmw+jNYon4bi4wSrBumskRTRo
YAwxPmdDyLCcoQpT9j3/x9/PVHjhibLVjIPyShkiuB81k+giAjoNEJm5wLFT2Ko9Y3GmHn8Rw9v1
WX8Dn7ITFpFtkL5H8dytChJuZXJGd4TKfnD1zQfV4IhTBDUdEsFc+ZC0Sy2FnEe6IybWMEZ+3iHB
supczohVy8wT04RxYyahL+1XYLdemk39J1xiUtojdmfwteBCvferL2ZeJfEQltY6tyKyRdsBqjw6
mKnoDMsGJ2f8imA9alwh3GNW8efn2MS5CbliIB3NuVkEwgGju5NeAkIjN1tCTXYmkWMk5oNM2xGi
AuJObz368/E0J9VBIdMq7WVgTEqX9UDCdfTMMgCQiEaomphVfUK+7lFyrelLCY7tp/PZroVjq1Ht
OuUI4Q/zjrjysyhLpt4w3ivWczcPcgbWZ+CxkmjLbX3R6BVdl/l9/uwkFylkoGPMkV0hlD7wZsqP
MiRGKWnSUSgfdrRTmC3ccCiIo82nXEhCIGHRK802W5fMBsn0iNDXV7JuFFFBO3ZpU8mtmk2uMJBd
HaO9RKye226SUG1ZjAOTKsi84VjlKvuJd4QMwTbmT0mUROKB0/IV6WhPMs7luIsmtk0koeC3BXcE
dCmpqKlYF/zhSTONT2UQCt10qL6ymygmQMHhIBAwoWB4vkinPrELSQUVyPzHgc751/MXUe3juwKB
11PTiNhiPRnFDVP82/pmp2rawfJWKpMz66CK5r6Ml2uMACQmU2etB37d6EdnVYXklW7KgQ0JICfA
rtW4rT4SepG1igl1iH1bBherBaeSRuGPZ5dN3KVlHp4gQyjTfPkxvUdxp6gHK7eLSFHPD1OgG4Ew
JxtUkQewB1m2g95SA92f553dymBqoY3StIxccW9VSBPopDxY+4jDcBG2jkYnZtur3NR4sqnAuA9l
sZ64uAhy2JU4YUUHTRIYglsd7IjBvM1mq9/FaZnJ4/73xNeb5Q4qYUGVP7jvzx7Et31bvCbASRz9
pk5DfIvHEU6f13BCLEmMik6OGINOoVdAHEkvZMqGr5P4dstQoPcdsxxS/KtelwJTGODSy9BNrW2g
yOBuJ7K56Sk7Ee5Hq7kLAzFfzMDq8WrDKGDm9ShaWeuPNEqABcI21PBCTqfpLuPjXJ4/nsAijHZd
c+6QI6mktZxz7f9k2IGSHV5SqTp+Z9GuI+wcXAtwxyZaza++OuYj9mBr7qtixYOJ5tQnsmTes7xL
8JJPY1f9d+vorwPsS+4/pchvxtk/xmCcSSrK6eI0RLC8XbF09ASb0QcNpowxBlDkYcWX5bF2JIBW
soZ2T3ktsNc2UOGW++iMhBc8arIc24pUFoAkBHgsay61vgN1a5pUSUlUdxtqFW48AFJ5R64i4aZ9
/bwB+gnmhlV0akioEw8noOLeViGVjF4wpXgSBbxr8TP52TZX/9xLSMBEq0OO2HLLbZa9JmBkjfcA
cIYdHAXt59iRQuIRKqUdL+c8NX1m/tCiqhHOTNFV0BVqOAwOS95odSFK2DzuqA1FM59UmvxIwfZ+
cBdVzL9CvDwE6KJ0CC0/YxO9cAP6PmG4lP4+3ZtI+8/TKVbm7y6cCaaHExEP+Bb9U+S+SpdTeDUF
vsScyyJebwZdRZyW6WS5KWKLa+6WwwSy0MpPB6DeGSASV/xkjOsURY+xs5cZIZ5RkkD3JXGyWU30
69eHsIXMVcSZxXoik/x8Ua5RoniDqT49Y51W6NmHIoJ3WrKfgDfEdwrKaGocifrq1XiH0zA0oQuq
KBpo1ISnUCUt5rNcwEd6LIn1zeTJBaq6sj5ZboOjD4SwY9chvDjkNzzfX9zTtqXdsE/ADnk5ZzEs
J4EkRj0493+pcnIukWALGDdHok3bse+soacXdTvnRiRVWF49dvmdjeATIOUgi+CBl8s95ffRA6Ce
rthf+9Vz4dMtwNBhJl2kxG+/2I7UVZx+qPVL9SPBPnOTcJ9LNNcpGVUgREygoPnMgmuFUHZ54OaM
r4tbYIeX1jwXrBK8OFoDMbMoRpUKljbnl17ktCir84qI/+IWajDTLEoJBrWmM6QsCzfiMVNbiXBi
B9SBzi1Ly8uMP+8FtdsA6VX+ERjJf/UXSCswEP9kEqFOQcY8vMcDppIpK2I7MFjLkVYjzpvWyF4S
u0pfn8v9Nl+LF5mz3pnMsTPGJWvUJurRlqqx2ZBwcR72VGgiJZRNjxxKaaeNL8DussS9o+t2Oey/
IuqM0Np5QgmWvZadIBQ6hliKEloN+/jfEzEUkc6qBXWJWu4NNGnC8IMCnghVtegGZ9fXNnpsVs4V
4D2MnpNNrZxBJ5oE4VDE23w+/5AjW+MwioPA2LeOUhFNKUFtLD6EPAdSkGWEi4Wt8joWPF9O8aJY
ZiLG9Y232h5AH9v5EiAjAZGt9Ig9j7UdlBwTo13RRQwwtN9mcywnp0hN7YXUxPWNZvGgKWJ5ROAi
aGRCHiqTxQPi4lOlwS0E98k9Su1ItdyaM81a3TVFf36JNbMrU8SdASuxfUbH2UhPTt1zOpQ/zdLx
yVywH64og8t5pZtcqLwuPqgRI8sCl5cHZF44QjgWFOPo8cxssS2kcj3D7xuuzjd143gCYNN4GfSs
dPcHJ7c3TAaC9oUtCnVhkTUJR8ARlwANuxf1U12JP4TuihVg8Xm29JnoW3IZgrHF0yQUl1pzbat7
8fE46X33fabKQ4iEc/CB5e7M7dcIxnVBn2V8cdfmhkH2WaPPU2pA6ZJltyEtwmuHz57+xJURmuqP
KlRhN7/yWBiP0UWBFAavVxI0i1DHDtxplfYuqeLA/PUl/EVBfdXI8oonfGwwccJ2kAkqrvP5xR9f
xK0dfesWPDnctHBaxSUQdTzACWSNaggcPANM6iQi7uSM16z8hjGJIepPRM3Ozudgux2YwvBLeJpk
AIiBsJa1FMztsfDJLdyidFh+cY02HNScqir1Zf67Vie4jmNIuptrKSFFD+o+5VEDg/BOkjGW/Gzl
ubDw3vVAS7ItC15QZ/AzbiNJF+dCodDMDEG3WD3/Vgx85gRsvRA890ti7jfVp677shkpv4p0ZxOv
9hiNoOout+R7EI5flyVH7BBN+YrvmzC2Hwrpp9WD6tURU0nUincvccxl258eGBlxw1GStJt+n+9G
OJvEPwcRdPPYUqJjC/hM+F15c6CcaVSkc1FpFEE0WOK0uiM2kklFxXcY0Ne9mNL7kz6qEqKZVHXa
N0/BioE/N8vNd7sQIJ5UM/6lmUINNlNJeDnW6kwzykaazDFR43D7m/cJ1tf8OsDVgqTq2G4tS0qy
5wKxmab6w9itbXgi8v/vHv0kRJK4okgwLXub7djN9l0JmtuotIoxmw1xKw63LfxbuG9HJgw4wdL0
4Erl+QI7LEwzcfq39HHsotcDj8lExiqhkUc2FagiJZWcyBbAxfqHCZsLU2BVD4J9nFEo9OwnptYS
XLNCfNtNvM5kZ5leaTjov25ZRht5fnsIZ6LoH+jb4952YGxWuPOJQC5u1Ew7CRiq90qpFi9VPB40
dro03Ig1FSsPyInZ7uUawCYqyqioJMPXIA7iAqAxKTrHAONxQfbWusp6wnMph6JWS5HsnaNz/nU3
eQyDl9ysnaR47KgEaDOU2ZctnKh1vqVhlEX1tEt3NS6rtmFW3oOBcDSht5yY4HQuR/AXsVF+toOD
RJgBlf0yM8B27LaU9cuwnYDsv2x3DmTY+t2AMcVe3/CPRu+ZbafHVkxDZ4muAlc37iWoH01hWJl7
n18J7m7vy1pdhh05Pf9gEjizX9zOlSgY1E+7fJmRSftKu+Y+S7NukQumOx6fWAf5eYj9wqnLmpS9
3Jv+CtUrf6z/SSI/BM96KWGVt9FRm78LjukKCCNl3p6K9GO57UOJQ4YZn7DbH15v8rbWgHYzoGse
Ix4gn//vRJZr4ngd+z5ASx9sbGEZsIrzjB8LDAjLKA/vSORkoETNlV3rna2w+JLNvE0s6xW0Uv4C
+VBsX/vOn1sU3Fjc2B7Yo6k0yUSUBWSddqCuFmtj7VEi7n9bnfAorpg3bYTQhGOCtjwmtwgZErrf
gSyJZukLGWGAMCkIH3WBnu++AV4wcKhEocMguSJT6YZdjgzhQ2WruZBp7xDqPdwXTeHu7vOS4cED
5p+v/Hul3trjxMaR0uTvS2ALvhOGsTVlRe1R+Vr1RtA1+eNbuJfSBMEcpC+Zd5t48AeFuAogjHMQ
d0VRkT31BsZBCPwZ1SH8W36apNNYudgzkLgoPS/2/npMRfoDkQnQSmnZ5ja/m/J3mDcLGSVMiJmj
7OBNwN3o6Ur6+VFKoXxPs4cAaXpPMSdBcVRSLgSxmKoMKJy70Rb7YAmHPHSLohhw0wsD2lnhhI7U
no4H1S7VbZCQvxJp+lxXvKrCqugbpRwRhPZh620EbwVQth4XsnVnp1BYpXXkXb8nXoCcY3+srmir
2hs8W5IyeMQOiVnGIGSW9a4ps4jpoMn30gdM5L9aRZrfRuM4AJWixV4KvzA1v7qYpvwfgjyMYn6p
G4P15ZQWl8YtZR8u42ES8nZ+Qjjk9uo2MsyYtAdJ2NyUDW7vWPewx1PdZ1SjrKCEvpE7RzGlFGC2
Z8fplXmxhelip6poGCdsQlkThlLuJdIzxe69ZgXDM7Ro7e5yED674QHggtfcdb2sAZKglOntdVPN
/9zrCZXsgVXctdEblZSu2BqRyM6FPiOK4dAEf6RtWwV4zpaL+TCqGLHiJpHs36Ys8+aBv392nP7r
SG/eD82O5ZsHHjdHZG/R8/PVH8xCqkZOHCPHHWHqt+rh9IoQQ+ia6vG5zKQQ7yf6/XlRiiul61pz
c0Z4R1OluX5HeQ67ck1Mpgo1PmcTaphKuddL+BZRtFecoqdVFrnupxrI2I+iHfNUCdPEdPZHiPNB
F/bo66aY9dyLiHX6+Ph2kWM0lPfZQEFQtu32udDyjdbzUTGdAKk3B2uc6e+wRXwoReGtl5Kzuwhq
yLUJ4enKhpDc7TltiKzhSUcHgX6KncEsl4Nyz27koW2zL8g5FpAHhcROgyBHWcUbFnAJCtiU4iUf
Q2p6zuaLM3vB7kdn9R9V00k96aGCxSTR6JxFCiY6BwkRZStdCmVNoMVooHsXbeGgGIJ7Om15MuKH
jUZ+W2kdAWQCSVG8I7V4rajfSvYX+HZPUMa4OtNjFacI0Os8Asl8fOpQWxP5fcFk2d6KICO4rH3B
Oztb952FfyobW66r6OO563N0oJYdiJXU9grTrJ91QImZbCjlBT9zIEr4eWm7iCPhKpMB+XWKoYee
n1YZmPybMK+KNr5M5srJ3tPiFlF3ZMNebccUus1ElN1LmpFiDjLQ1nkRJ3LBdEnFzu+l1XJ9qrfB
HR6aMHj2ZGDE8y+oewjjtmamyObuBvdWW5tQCNQGkUNfF5nwBxoRrlvCvVzFPvESBgBHHONNGlx+
uAgtxQkTSg3+hg5tZQtCN180PxmBWY/S21KwKGaNUaNFjiW9naKPCwwzJ0aK5cSFTlB/N1NfmSNl
W6z1uM5562lJAuqIEc8zntIxcPCTNAa3HfdFcV4AWUJIlgmp0xerEcLQXAQUvRSwuYrlJmcJqzHh
xZ9IJlkyPHcF5Yr7aSl65rS3Oj2G/DBeovmiOI0UcHpe7NrWd8BWe7ytkRdN9i9hQgHC0F945kH3
XL4wf/yFqmtjsbiEIoJviBh5cSY5imecjcQzN7b2d677mdFh0P0kqW3i7tboOvmWOzEUjU4C2ETI
ckL7CW4vwwd1uH9V3vSPASHJGGJVN/BZ5g9N1cxnU/spmgnLGulq8LY2zwHV3ZFLB4c2YibK5lvq
19peq9yod6c38DopNpsVaQgP0Zg3MCqSLCE3uvk6bntj0SHu7uPogHZBZ8+Bx3c2wD5hweFabE2l
3LR4ppiFn5B8S65sr1ScicZcwD0yetHr7dCFgszX9sDXiOKDscfm+wjd628ZvRzPNzyCRY6xNqFf
raYYlkdP1oKpSPowtaw5lU/p2NO18q3ar4HZuq7kR2My8PoagaQMaryTO02uvH5p87zU89kK1vTu
uEI/k1kSpqkN12ovGyLhOCeByLwZupqKRsj5Q3XLwuYaM70/bX17GOh2D0NkobFeOIlhDQyO+RZJ
CD2CZ2C3zQ4REMRHG6x36iNaAXe1fHPkbXNzdsqa3PFO2UXQQmbmA2RqPEcYreHU3ay7XeX/xXQ2
5xzLS1NMy3SSHz0gib8uGd3skJ/2kIve2i2L/qC0JgvUgMYpch1gtc6NXzz683J8c3nPDo9QGK3z
mgu2T5ncWGx3sgJC9BCHJ7EvBe2UDmjhAkVaLpynKfdo2r20vWb+Wodq49Y5HkpDgK0bJDVSG1Fb
lrtLEEgp8xQI9ReA/PC3a5FsglelPtoQBmqy1VlZlt0dw9D7TU+FpXKuPmL3PgPvIamxJb2VOrgr
Sot65OhF8O6dBXo/sasni/RdQpMcge7LBOD8UcPMNv36V0wK8nZ7u3KRDHFxAeTA5Tk7894WuVMM
1FpubXt8qK0JSqWvsJ1syKEx7dBMseKilaM9iNteytuHAD6fJzP+xDIh1ZgoNZNKMLkocKmpST4Q
9iDjtVECybUoYEhwdJootLBcJNquL0FWPbLyFRbaFDPsDDzOIg3SCTestmvu9bvzJvno6xgSWaSb
kLCDPaCkyxXHZOzrwJlT4i3M6q6zAHoHHl61OMcCzBno3/XlrC6Y23vvC9/MSxl6fgPksO/Vc5my
FHTGnWfNWLNp5acDN6I7q1WuXPwkwHEbqC4lJ+D4RMkCcrTeG52e0JTa6x+O/uEL95bvB5YvFL54
EeY4xLs37YXk7aSUuTW3ep39ZD7oTWs1NY3Xnf9wK5XJewIcRmj1x4LGaPaUJ7+eSQWOWCiGAX/m
icVQ7htKNIe1ftLBj2dNpQKPp8ygoedjQ9uErrSrV7+d380AGHsAAeOu8qs9YMhXZzuiQIAI6jes
+sHG80MAyD2skVaqkTJAp5gQIoqkRJVNGd4J8+1/wrf4yEhdeNkgVVVYUpsEE4BP0ozA2KCBXdwp
ubuta9oR0K+yHXUyzav+LU2fFpS0yHroQ7eDccXvhj6bT4l8aZqK4yt+vpHV+sQzdtsuALsQqCgd
RLjh9fnTn8IMfyuAcut7cGHJlP72Ruwissv7CxoKLlcNV9lbNnFc4iS7G7q6gRGw2tZ4QAEWO6O3
u2E7M8wq3nrIidNt8VYgod04rtyXBospg4EsUNu4mxQYEhS5oh5URcYEGEtBs1RC3DQr1On4yrPB
aHr4jKIMFdILcYX2Ieof1V1CokkrcQPN0tGhPyrum9ts92RX8SoZP1HrEJmhFygFYnjSV4evVWLN
QA3Ni1h+YUvxiLoHud5CjiA2o7tUZ26d04hB7WouIziUthUsnBIV8KRf4qxrprinkawlQKOKNMjD
5SZjhJ08HrUxh+T2V2shWsR/d08d3i8PvZ/qErsO1c+GJ9vASOKKUPoKKSYW/3FYieloyUF4/TXd
x55TJonEDEUmRNbWH5FWkYC2Vv7M7t0i0DsDn7pMAfTiv6uJsh4CkU0w7FBWI19C9uIXH/9KbTOH
q+gO5/WCu8lSiktGEJv/2I2hDVBtejrI5O9uzlbBd+yIrLMtsiGwRG/7qj+1gXy0f0MRqavY7shw
3l6uyCutT17dVnEqKAmqlPJG7/RGHQL/YDZLMmiirc8YsVR8r26zeNL6mQxnLOCAoGTfMFnZ+shh
5HzkkVEuf7DBTuVx2cHZzk2nYvqutHuQAK4q83elOIET9aG52Z6JUacYXDyQeMzo2c3JBDSR6smm
vysZQiyix90ga2yhayYNLjk/jk2eSSNmdZ0zC/6WN3aj3KU6w1eBW462B2T39MpjSjQBdJv9rvH3
RDthXSWVn1fCOLEkAp4KVOb4GQ6gm8tMNMgGgubs4RUxhLY3A+LS3LXvB93ivJi/fyByGLOAFwQ5
qd1xWKqLarhU/J5i9E8ISB7U1JacQZvA4Houw2xFWkRKGupMVmPcC2gh2frJLX/M9ev4zhJUfF63
zCHHLXcte7LPxD5bkHgSBz/Pr3o2h3LNz5f2hn+Ykr9huz4ou6pozyAA9shLnCnStnBMS7L6FnIS
JS71KQWViTWfNfuNJ+AeDdMxRZLArhSdEAIMGYvW/VSt4bMzevMdWNl3uzvv3i5hImrBm1mdXKap
AfXsLkMGl6sK+dfNIeXajcpS287wVPV/SdbKJWRLZfLZ7bTFoiFIRiZnvBfvQjbm9YkZ0iChWrlB
DK5CojAvYdMALPvTBkpsiGntpu0aiMgAP8YnVA5zyzqnsmiW2LpFne1+9tthLgrV/CuMQKI7qiw6
aJllrwt6AopklYW38zS5IfR+317URuduCeTfEzaHrMPk47tKon0wNjiv4/h2yi/L1ekzmbBL8NHB
T1Cp+74YvQOxd23gd/qfWTTemnyZ8d3OAjJe5WZmX1KE4qcKrQOwkMZF3yr719gJbNHpGAr/SVBR
DHq17MWQ76emtcTuKuep5XNhO2O+XbQgAs9YdGhGAY0+wF10QE77YTrRNUoW5T+os+GAnqEBqPzc
DR4kBDPkMWn24QAbZ6wnAuTOh+PnICaBElh7PXGYkGe3L3Xak+LZw02S2FK6wWTpSHOTWqZ+5hPF
VF3vMFfX9G2wAh8rSqgigYMiLbDrsIQ3FvAgP2xjOt8Bi423VgIqoByzJ5R1mbJg4lUZ9KCBPc5d
FsPtD/P0rthYp2DSiG5nGaOuf+zRQbF11HHBipuZw0gs1gqnKsWOscuE027BuS3BXWCb81UOyy1m
SfK+SCJ5+Qle1UqFRx7sg0qmk0uHf0OaAPsIXRw7QOLvCOgqcWp9417U/VF1MN455bWpsmFS+h0w
cOkJfzXc2TOjv/xY8KQZDe9Jmjm7cIxIlyE35LLZacMnsxsnzcPM7gnVFSOXtsxFiYiVGVxqg9lZ
RyRWjhVm5gRz+2ymDCNeaFAkhrdipfOsRh+mdRhvoe4k2fbPQAiHGRlAngbt0OgnA9OyLoElX42t
gAlBmXty9Dti0HRj345+F7iED5g2/lFICBSB0aPGf96uo6eORgfuMhfQ/OeRXuKMmuUGO0NiiOt5
H3JFQfhCuJxROlDW8YqnisWSwlfBgUU42meKxjE+e6L4UI8p59jYQIkUFSDDq+VcOYiT2pbL5ZWW
8jYjAW+4+BH/V38a2++vTdioVuVYQGad/aH2e2BqHyoNhbg1l6ybPtK9BNeZ2kzdfhPdTutIvYp7
3yQ4Sc6WrL4EYpfAtwVMtwlSlt7Z9Ef16V5xKQ3LErBuYa9fQzwSpZPHW1vJ0/eJat/ps8PV44Gn
Y0Qj3MgWnLfnsEyCyllK8S6ahWfOIy0ySyvkGF9k5jaCPrQtCvZFITfk35+CYZtVz++WL3gdAZL2
pd307EWjfY0BlaKm8/Bb2l8OFbjpxjV8ESTpxrkE3B3K1l4egNeas1F/s5T+bXLAbUw/SskiZUDG
GrbaAaWlfKqFOf8Ji3ovc2jRxD/S7IxCq4uT+1L5O/Y6v+VsU5PL2iNwzG6SJLTif85p34jw9p+k
y5kQICGUgk1YabqcEDQpczJklobnHSqdrVbWkKLBNgJXcY0eZtaPWcOFNne8UUyNEcxG8nP3AZPa
NPdJR9nvLfQPt3nsdNq+WYXh97xAZUq15SsL7JCIVuPuU/3AVylTcaKKk3xWEPYwODbnsFnIT2K8
s8ciiFl6hj8duerdQxHNMKEC7m+/jYNEF6bwClRQRkXLH45AKZewyd0selJPfNKmYrq3A+yFrkLH
ptfHtbKQwroujErO4m/nkH55tMrAMVyz/VD19UHDxP0gp3Tdm3puWcOcyau2ktRlxmy13lBEdZB1
Byss37k8gqLXuBc6sGlcwgUsv9/tFG/T5Qm4AKg6Itr52Jkni8cJCq5Iy2EA4rkdzF88J/3ZYD7a
6u3BJrAok6lIOXPMikIQa6UYLYhx7WSsmucjwWO0Kp7lTvYGpEIfUNPstskh5LUDvaPLhyoU5ewu
F2jCKM/OblVAO3f0uAczOZ/dg7krqCgvt5+zzGOTUUr4UzwfrF9+5hmmpeFju7473c5fpti4+Ib2
HMheGrHrLlx6UvW+GObW+OtfAJrcVcu2Fz2s9PDd81Wk/I5a0CJRgF8p3MTVV45wBZxkPRllRgIW
wKkBPHnYAJyDpg5sBLWt9XaV353ItvABAMY5OfiKz772zRt4RUSlab4cYr/6Buhex+VTI7UwU751
WjSWjt2FcReUxCBu3dC2lLj1PmMrtdCXQuNSmIQ+hooh0f3ciD6XfYQK9o4tqmcY96vCOKBX4d40
3amKfcAWEyGT/GpU3b1S48VW2DUDsSQ3QkbhlqbdK4SR+CWhFnMTN1LfFVLGNbcFJxh1jN81J6CU
WB1fbhWAQPrRGYBzrPcOlFg5HngCBcJFzLLdvPpGv7rl+G5A8EHvr75wA2dzyFew2qpLuguIp2BO
t8CP/p1Xny3DYKr5SFB8fplHG49hDhlbrpGr56nYGYrAM6cYWnClWP1tDQ/orfczQpq5P7Z4m2gC
MCf4mEFwWxwCQjWAqDz1c3z9wXRcJnRRjmtJ/kG0hmGMKFvnEv2hkTrSkWVAUNyCpV1tmCywdYyx
7cgIZHzNFWImj/p/UnrLWuggS6uEfuxmR0pZm54UrBVQUr5KVlnrqmpZ3UXMRwWxmwqusYBgcf3O
91QJ4mQa3VZCenwqlAW1Uz96nnJWTBlZy28K37bGiMuzwyg97zBOQ0/XNpoR7PsQC12rNnDu4vXQ
4mn6gwQ9rFVzuyFcaUapINH4ZSl+rK8bMyChV/aWBUos3EHiVwpp9gQYzy1LJnVAqwTmP2hVHwdF
TqHNF6wncEIDC6n9cIrpnnYHl4JsQKyR5hNkYYoKn6Eq9OUyTFzQtLlqbQ8CtKA/VAmkSiKXqUg6
iznxsJvQZx8upHS8+NEwwv8ftzesoorDu3918RCWfW3LTDWpJ1UBkva290FbK6pT81Kf8K1Dj+3N
eVk7UweOPcqzS9BCYQmrxTtAzfSKLPJZfwkm86yqMbXrR6ldjzpIjBmtrJ6EezOLE/SO12kgo14h
kDFXD07Dx8hu9etH/axJrtFcsPodQeqB5iAv8MqoLiSnSsHxqx0fzPWMngPr1LWRbTY1S+9wgxAc
2jg1kezHJngPrVbmhdb4gdakFY8lMiudxV2LSvAFuYDrS/9eXkhEsIODcSyG/I3Qf5O5bhdCxj2O
XTnwENsvB4/q0ukJc3p84UGITX8K8GoiVtfT9dB8nLiJUicGo1TbGbtI5jEYl9Hv/GyAlOCNCWr8
TUz442unKHyeY5XdsWMIAGNmvL9Xum5nn0iVQSuH1aCiwZc7HryZab10UcIdiS93grU2gnYo20UU
IfdF14jreo6vxR5SHG5MHGixDGZ+DsWTheFTmXSaCv2aUSt6Ua+fWrcvsrDGX5Afi2gVRbpR+gee
avn1pTLg5ihI2wpT7l9TuGGOSP3nliV5VgrdgUgKEgF2AACxHDEkMt5ByZdc2eJdG+7LrWn2/1gT
UEaBFZ1qV57tVgedGfoTKrx7Mbc9YyAQdIDC0eFOi8UOM59hru7KFOhauT/bvxsigxGlY2/ruj96
bnKikFYzyU90H8/Po0h5LRbeWHlXbeNQd6sVagH3mGVOcY7WlJHnyZMNW68iOqE8GpLJl0jVbH5n
S15uQ6me5U/54WPltwhaMVh1wPEJtf80/y9xYUWQj6IdP1mXm8PAtISJGFULL6BNWEpm9HupUBUk
rlvC2gr0esdKYISWa4dulnpyZdom9nsvzy9J9NFd18sjqudCvn7qEILl0v4mh6PC/WAv6t/L3Fth
30+s0q2C4pjpTXDJc/7jOcvVKYgQwuQElDzjwY4NXX2K/aXKm8OKuyIHQlhsWXA5gnp5uZQDTbgC
aFHzD0kjTI+ZgyHconENTvcu1LQYOkh7vB4EQdLFElO0JnJwEKjypfItE3s/Wv9hPhBBdElQkKT8
MUNcrDEZsTwjw/dCFhCLpcqKREIBVDtFTUGoBZBRRy1zFFZWUICqunv7dWy7NuznqA9jSHpEVqIX
sflulj0Xq1WSO3thG7g6wQB3pMZ4n31vVDOMKSYHx1HGAf4yDEHM0g4nKJsUzUIfImuQ/ARlL0V9
ji6ly8ZcQeFKaU7KDgX+pSbr+KmOvyJNR/t1VTs8bVfgcdw7dEBWeRRr+13Q2WFfMng0OQKCmCRs
HI/uy+24DOSIYvLLi5AaQ7oJ1yYqucfa3E/h3pyLAPvrKqF28897/jcxTjoa41EtY+4Q9pY8mxtP
jDj9DY7RKyCJxq0uSZYLqm+4GTM2v42hSHH1CNoxg1K0X+yGoB8zYpmQTAMOiC0j/wXfLwfQ5eyd
bh5HWvkbxrArbgCve0RWya5do1WMEO4tlZ9O4LwpVW++2igtX4BX/6HTJPtsy0Qr4LzAqI1FBW29
Cc49oiuoqOmoWJJFfvHeb0ebTlrIiOUUhCILAtEh9KsoOyFBfZtdnNGLuzivGJT7iII+KOZj8gyI
McK8uNGfJFGVxG6wpVpoRPHWzdAY7iVzsYw4TWg8aopbfX7DH273x4WZk4dngNkyzJsflBmSbs8Y
66Ua2Uab4M3sSr1n5kzhaKL9wo2oSMs5XfAP/2NZO0jXIsI1zrM/PNyNJgyxxbCcyw7vt4hOVutl
td0EoqxJACR+o4T0Eox587q13tifINeHhR1hvlFFwbqNvuHQhMZMiL984Wr+PcBWcM0/Szisyaco
3LMJS5o38S3aUt6BSxzf6sKdXFrNBNsS2MwoyTN+ccy9mUu5yJE9asLJUgK5+JFEAniYGCPDpBfe
MqVsARgCeLgDfv0J/iEQl2epvpNg9bTYtQN15rZkGO8OTLrgEer5PSlEsAkZoxOuI6+5x8UJzgqW
aNIwKO9kMIFxsJ+gsGif57Q8YyfqfN9hUf0kNjb2PWmQrjseWQclRRqeYLmm5pIpt61M+BqRlKgw
u41/C71aMiKkxh6cqvWmExQEHKLr+BFFp6R6ploHnhzn8jNHYSbKdSZrEOof8tsuErmf4MqYyfgf
AUuK/xhdFEE9yjgpGk42yvj4kizgyyJ0L9cOKXvyJM3AC0XCSHAZPLylhtzCJ41r2aqREFZfpr8A
bGvLPjlAX7IzndIS50A3hbmZbTlsfiO6mL7LFh9l4xUvvUsT9f+Tbm0sQb+G4ydYTbsgMinyoXXw
W9fGeom8XeRaKU/l6wnp7iGfaZNR9g3NFGYMkFyyiJN7MNDokt9KVR2VhR/vGsNMeRTPgM8AZUWT
h/XmgIEMAQ5ACLFcnADKpViZDlhPKA5zZRqlRAtPV6cIYssOuR/EhLr83yzg6j6AlG4fc2p7/OFl
OF7iEML/3P8tqBm838fldkShC5PZr1LfuGrIoGY/N/8aLxF4I7x6FJXh9CgzkfCnZgdWC1ARYW/u
9ZLssDpmta4UhN9q4vJGpI/xZ/f2/kFeHYcgmJf+dTkjgJwrhqdPpQTdcGB+l58j1jz9aKgZPRxe
OQE1eYPy0hBzMN26piZI+WRyvG5Qt3PhacSuM/HjnaSdI7UjsX7rLqzyGcNCM0z0KZcBc/zID0QQ
HTGDNXJ1baqtAS6V+hYAaO/GWHabautyKtHWMbIM0oMlYAQnKrVCN9dZ5clecXkMY0NvVSDry+kb
B1CAuPaaheCpCYN2l3joBMsa5VjMZNOK6BWTVKRPuY0U+Ntu0xDAmBIZe06WSoISX/teobE33Aiq
l6kiBJlkNnVJRcBZuSd3l6UzCjjINvH3/bzC669IF+RtFRfd17J9YwlnG7+4aTePmYss8Bh78ddJ
qcp459E1VLNTqlDPtxcxO6KQHzlObztwufmIspOQ2aPRh+wSJbTKQPhqPaDU92aV/kMxFy4Nd0uX
m1b0nYc5GhbRtRKmIkXCt5Ml//DvzOV5BrjbW2iO1Gy+smMnQf60CPVRT4c2WBl+gWwIS9RjGTCC
xhZyZelzfCi4ORDS3rOFEk7leBq+Di9MP7aOSEMR7ZMa+Fc17Uu6a6JPRPoXy4QKq4AgVIsPL64W
YLq1zBD9O3BuPABK6+kj5gLa6LGjul39CQNKzdCjTBPsjzBgI+PaxMjBYibLruXP8P/JLI0hj45g
y4kD5ceusOjwPWaDajCpNttcMdGwJ8OzSsaKhfduQeuFGtrUDiMICjL2p+7t2AWr2zC7rYXysTLB
VWrgH9w8GgP7W8ht2U3Zu+tX/GHYW+6v/qSdhfwr9XKaxmUvMsLWcIj43yB/pbnB7Z3U5YVQa+wA
BoUBCtva7+t37Edw1fXMLpAAK0PUJhxWK7ejk9SIsM0OXNOdW57xJPulaSqywnbBibCwpzI9E6b+
bu7gdRbTqeqcau7Zkedy7qq6+XX7qbvYn70M1DOds1GDEo/+wex9m/KrV6BxKcXTeQ9MgcHClkyw
6bty7iAAeVv4jLk41obdb37x6k7kRMusJvXU+AJ1bGWbFckp3WcZNfpF5Z+5M04VEsXuC7sdkP63
evhn76cdPgRY7X66JzH+7OTKMTFK1lFK1IMM8qxuRISY9acB0TVTmwzF38v8glyMWXx/d9VCKHg/
reiyDw9f3u9/r0GD9f06+wah01NHljHbFKe1FvWeY8U1/2HBoLpxZtAEk6K+VK5nJcVAy1xuU2pV
SB9mALivFXmrs1Q/MZ6cwuBVRsqo7MnkP6sUnCojnMSYr/TgO93RbyKFjcCgwSKx+KvzYPxq2Cn4
8JSJzEhz9ZNVqMXTrt5ZtM7bPAS1KYaPHTSLPA+9aZVMsi+aMY/B4wdYIERaieuziaR8IS6Y7Ji8
fbD5V0pdVK0LbU37T/34qKkcOeWmYJFpX+FyKs253uEU99lUsOZ81AryOLNDIsSSBcrYj66kXAkh
EZhocAJIpM3tClT5O50hWPGMrVHeHCwQFIdyFokELZ4YcZ1kZyaBMGhZzP2yMAr51somw2IK76v+
pQ9H91cK+qsM6mBHlwjq9mlCN/j99N6/SqC9NHUrB4nESIgGG0HVo6SomK50FWAEafw5ts4FbafP
GOl4Xwfmxlstht4aV+IYZHy8WnDMOKuGzUI/4cYGRsObGbfog9u8qG3M7cnk7M34RV0PchxfMsIp
8X+BxEied92ac7vZTHdM897zs6efg9zm8QyBBFXZ+bfzbxS9rg7hDzlPLkXs1bcCU3PUafMgEUi1
mKFsfTsb14AZ0lAyeewWIkNjlD/x2M2x87+m+y4zGXNI5AR6Yt5fCet4cm+LbB8Ien0BycLvWVTo
eGRNdA+FiVHOL9WHERylRGD9eqQYPJXll9Igb/2lJUnlKkOm5y/1tgRgB80eIryDkG4iypeGL1M7
jHxK5JmHOqxtoow2CWwKSQE/jABK+k/2sbnv/NgG4ZekTkvcOjqKDAsZZkr2zrMTqqv0nytglCYp
gBxCuRXi+0l6j69Q+X/pcD0ESxGIc7LM7ETF/xjVt/Q35G3NGmoatdQhxWATbwf0ufZ4mgUZhqRN
bfUGDThqI6eGRvvKMSWiD0464c9WOVVA33b/Hk6+qOw3lHJK3OA4H/1k3qjE4vYD5MKogdRcnJ95
0k0qokRjq11YDIRqaMfpQoTdkDiQoEK9xoIEQqn5cvqYxu9tL2ohO8LXP0wPL7HGi7R3Gnuu1F9a
Y/sfFSbkjun/GFXpKAqwLue/8k57zi5SISjPrdjqH2wa+3GsiUOjR5y900EiYcxKrcRpOtQvByiB
CJQB2jnwujmw7LQK6e+EhckbBcV3S922tOIBWQTqfvc0Wzl4DF1cLccVqDMO6Q1eYSNZ5qwCbhx6
8NPhATTEHOp4pEg8mUiIkTrXw2UE9vB7b2sGv8ItvUWPdxcbSSWdlPDIA1yaC73LydbOE2IbRRWB
qrmzQmt+6YZ+azh3X59eqNr5tiyS45tI/R5DmwG6XOoyAXdRl+FEYP0iWc1zjGJGxCG1309v0xSu
LUh3aSLr2IGCoI28vxHOp8ZT1m9NX8x/QrPX0FVllO5a6GvVNVxabv8uKlzWQXgoYxnkugyTJ4WN
TZom807qLLATd/0PFknquw+IZYpSq/chVKy0LdemCti/jA7rtTFV2sllp4YXOTVLTcexu6zJ25Ab
Servl6b7Q7kTQHe0lqG+fIJdnRGKKJ2nq1ogcIFi78iYVXGF3Zjb+Iu/Pek5WrNO6JaZQLDo/xYZ
PjRASQZbEGEZ7s6u6ILWbDecP4UzH0lCfhl5rKNhlS6MPV1xh/xuJtyAdq0LR4XLLVBVdc/8XI7W
d8feomgYhRGHkA8KN3pzyaHjdXQxxCmIbWPN6bG97W56HHjRcxpaXM3MtU34ZBFi/Mjjx/tSYhZQ
c3WzNTZDGB2U1dQbUzlXsPcXxT+j+EIFbSrgg6GMJbjPNxcozMJff6UJX9SZkvDseDcXjigzEdVQ
Uv4cxt0/sgLh1uvSJwnsQmf/VG0gpiMbA2LDLobq9HM7NydZ+SMY9hdPcLLUPW3avLoAALt52Q06
vuIp7W4gXg5lZzd3B9x8x3uKz2bGf79g88m+B184yhmCt774vq7hYfsuHnfe5KrU0/WajJ/zKNco
zFwlffNcxqX8l2Byb9sAW7GGBa6+XxmS7ttm22HxzvxR4wU7qCniYnx1GWqOHX9Uu5pM2t+5onSo
7ShPCm6HsT5B0clXU9wIiKYU0Y1rIjZC4/nCrw8mGqxZ9P5+TCzAeIQfCm9NWIC1ZRpMtMTX5HLt
tGbt89DuBnk0tEEVa8KIPBXzaS3xf37kl/8GM/o8vFSqme1WmEanZkczkXHPx6MArTGi0vQ4Ot/0
gLRsKSLSUQZGqxMtRdkrOAHgofaGQcb1ZtOEIBuN1ew83o5F5XHulsHkiiIvmaaBUZYjZ+kuduQr
/Qb5sSb0nS59avL6OlQ4Hg7z9S6VelY+9PnCb+mrob1PHpooJjYEd6nblQTjcgZjRlM8UovfNxzx
KjAe6Dat/dWr3JMnshirugYVQGwrc0aLMnJZBHWWeCpbESMWzoRWUm6l3X5on47f6j/vnGlYU2/5
xlIxd2W/bMXTV9Kd10jecT26FXupZGEHx/zEvtJr65qRLRMjqkEjraitTi7bFrW6P/UCxSJngVl3
CljgmFvhahS5it5ERSwiuN44bCu2VHWHoAH6UfMei8Q4jVQR9tdSIZX632p3Vzc8qmFIpFVGz1xA
PtR8yapXIUvW6IKTqxgpBeFiwZqOIfEQbyNpUF9emc5ZUFa8ntTkh15tYlbAWzTYWUNwUA3k6tFc
YDDUXwTIQDoO0RwlGf+cffpEi9OkM83vnSDQzDwSWjGyO2l6JKFTnSLDMxo7OnIxC8sp+koea+nK
Uo4lcRLXTfVAL+ApukP6Rd0Qs3EEYSqyDv2TNy4FkbJlOUVIODg0YChgG1WVboX9sDciXBnolfF3
E97b+KtkME+dQ60mZCEEBeE8mlBx3rj3cvN817iDGYpd270Bt/RVahRMYCAGgiU3wbtkJ5kiQqx2
OEE/J8SkhTxb1gWzyScMc13NEKX0SJnsIjz2intZOSyDK1isK0tJcds85TbOMIUb5FJohcC4LR+8
vt60urg2X64/2AjX+/FoiDwHlz/WxVKk57jhjtwc86TNxDP59UHVmZ/NOmVn2mjpfXnIgAYJW5+c
jAFeZkgn6wrNbxK6gAEShE4kdXJ/RwFy+LiuH3UbMu3bEvTcJN2t49XdQpSoF51Quy8IrqKzMuJH
WV+v4Zb7w9wRDOQGjb7RGGkN3wUlxEpSh5zTPh6ZQzs/mXNp51Jah2ZrDeYNtt2IcX1l+IKp5H8T
oQUycMhgVlyCKimdmzaRF2lOVumLd9bvC9niQF1UqcZ9tdQfG1RislkBYIAfDze4HYOAilPsvhGu
T2+k6dd2upcM6EvYfKyk/02sEl/K5JE8AVnn7qCmO9VGxoqF05GKhyzhe1EhlMl0xTApNSRE018H
beDpJrtQnd94bi0raDWNt9QsvDOXIwOTR1gKPVRCWh3Swj0gmzjA1CB3lgYo54fH9y+GkmmbrjuO
6fBlk5+F2SBQxDAV88fIt8jFEoLMzFuZgcyf2iTaaQd/1Hx2ZTNLY/7kdFGZVJH8e3t8oCY4IzDJ
iB627Ayv4AKj0rl6AuRQ1n5GbfRnuon+/QkHPYjzMRAlInRnPYcRuxVxThXRiWS0osnioem9LD6N
C1KHOEHr60mrAeJAfd6gzUto53jveEtVhq5lyJ3HbCa5GpoD232e3swllnp0k6Sy4EjwIyMJMLNc
b5em78ZRYuD0/uHjpTDvpHkPX9DMyfYe3RKFapo0TN22FJuSgv0x2rpgLa76b0YyUH3cXHG0lXax
i+GHxxzJwLjkuB7IdA066gSXzwSTgS2gqgp5asFtcvRWRPtLB7PNwXXDpNAwxSINv+3iz+e+MfEK
GW6hgEHK1q5cgF1xJuLCf5b0o6MZv9zDcAvA58FI049a7xveFcJoyXrWxraVPxNYZ/+oCKtlvOup
TN+MTmrbHRp20+U98GZgFEBrqb726SLZcSI8EdSdFUymHYZt4XBv0asr29hBkopauHRllWkysXf4
+9UGjMRE8X24Zxs1ut4s7GUkLvUPFRTUNVlMA0Rfwt9IlURHEwR021YKl9/YzpuzAHfA7xqXxbny
Cckr0bCbrTfgyNsinCzxNsQYzU6YMraLsL4xTkQOz61G5p5TqYMwtk3lL9LHs3jOS3iyN+SUIGOr
QeRIIFPJE/9HHDGUEihuVRU3iViswRNb1vZ/I/uzm0HP5IOZSJZ8coLSz+JisxTqM4RknLfBRHNC
LJ/BuqLodG1dUE6kj2cuutOTW2OwE7Zi5yYsAzA20b9nakT/3gIiyiA/u6VLH7trXy710T8dX2M2
9PYJT8ByYW+/XpJU2sHQOSse+CqS95EGJmQ8x/ILlTX+jAnQaWosMLMu310m8LGbJ4r8kOHtbwQa
+n2CAwO7SJqacUq8e0jU+g95pGPhuA4xOfLwk+OBiV64mHMW4/Z2pdWFjlm790DZzKizU+QO9CQZ
pzickA4+mgrgIyzKaWUrZuXYb1pL7XwWgO69fH51sKBBSTFJfJ3xPB4vtXSXcx9o+dUdZ08o6bm+
Wf/lvQCLq4n0MZNdO0v8AQOsLrLokFB1Q5G2h6J+X7hh8Fscwxfhn0ptCRfVJrwsyx4w0lE9cMAL
Yu8Fq0mUdPhtG3V8SHrVjjpkPt6qlpqbhEvhEuDSaMrDoj6JHLqjoKgPHgpRmeKak5a3gVf9fQFD
HlaCbETFV5wZV0DdydOnGhVygn6oSRqdZBpfmofNCmYq/5JchLe97wwxgHcBNSr8v2csoLH43Ale
qMV55OC24BmuZXBAdu/bCrp1QuRLdQdELDmU73NG5tu045nVg7xXQsO9vC5Q7bqHQIVoFQNgnVua
Vfq6jMKkD4iBuD/8Z/8Rr1HVgefhk/1BGYSQVN9E5pfOPbJYGufE5N2QqOtGrdtmi5j9j4hLblpt
IRaDAW5WgOcaES2kh1Ksm/gseHJAWVxTU1jr86MD9taw3SIB3xUcv5IRhVl97chhOnwGuDRYv4MY
KO7cy1NjAXeZl/BoTYhyKyArYTeyX96ZeM/7lzrGijENdFWZq3D2Cu39177Q9uBRlRUE0WP0e1XU
I0l2HHToBRe5mjFiv94Di2fYTsWNid62cdauthpoyk+bSglDIPJUsGUhNabZBXXA56E7yD+jEzy+
6XO7KqlunO+aRrWeB2ZDa89nqaoJfBevtAmq+VdzVewFBs7Iqd77dTNlaEMWfyB1bDeRuEW1Z9xv
v3R+vnq1T586xbfEPischTpdRslxf+2FkAiOuz0mbfaCL1Ar6ZcvlOEf8zFrA5mkjY8JegnxyJ6t
oRREnpL2Rm4uwT45EPPdr2Ppz09b4eEqOKLazuq+mjyr5+59odPwwHkeDbBAon7kJ9x6r/exOBdi
Iaphk82GcEmqKXMmJUQQb7EsIaHpI/PyFfNwAuNRFR7wd3oERtd7UxaIxvM2XKq66wlQuKdmr/lu
EbhTenMaEmEE6cKKl3x5uVQY1EZgUDI87CRyWwVfAcf9//5C1PWXV/6aqH5OXMzNEH8SiEItUth7
1Yxfz297UgQMQOdU7HYPz4Iogzo7nrv11uUUh2CBGPSz5oZ8/CmDuO/BKtRsgDabH3uOvqiDqkou
KIswtF4e1KNTp7EuzYj/xoJkKxbmHrPifj88sIzRUqbUSL8BuOF67TWyJvWQ1Qt5rpUFf9T1S3I6
Piw/wy3KEIKMd/o8VFpveZLOU3YBn1kesL1w1zB8X35uSY+s2WEXcfg8edd0uWAqh0eMJC/A5yFD
Q5tpBrnhxtIJccbt1dhctyQXrSDTHYV6lM4UhSramv8JeIZeVPMYi9FO2rWUPQ7mdrXzIGquC/OS
/jT8z6XJ5oSiARyONgG/DH9K7iassRHLMyT4QUwY7TD/08qjYiSg+LgcBNTuXba0tDj6Sto/34jR
zY0yfGLUi0NRNY9d6ZX30kIv3+R2/BQt2B5Q7HFDzIpry9czK4tGewdCjJKlp6VFm/kSTOlkrGiy
xyG9nVyxhkg9aA/CanawEocyUQ7aGho4c9qNNwAC2bdNYAtVut8pL4aJ/LSgQFKpJfAfYsTegcEG
Dp77DSTdxZCjtkofRye1l+BWtXhjINxe/y2Jygz5UKaxKAKC55w96ha6YNmeDgA0/Ye55dMYjtwa
riOFmekWm61xCuulaFzMIKqbfCnjEdAnixD48MH6UK+VM4IFVmaCbgPER6xYANpeJbWIelGQ7X05
qM8hYN2qi+esPNOdYSCA8atKvOXE8wWokdaWp4b+x38B7bt7mXfB3qC3rRMC7jYd8ROVCegKxX6T
Nc0aO5OjM04tgC++Zq/TekS7oYTzH067wr+pjDNLlkOM+0bZ5f2t8U9JbM6Y2rOn/UA1tBQIJBZA
pmy/DOsHFFvVe5uOGked63iUCN3dTUV6NQMMkyeE9xG6yaHoocAJg9pzUMqbFqeXjViCdLu5b9zu
TattbxD2yPeD1Rz32za0UdGUV7IKwFhA5qNNl13DRmCWTJaBrJS3uFZ1Po1H8aG9oSAnNTiYVucE
EyTFVI3C0Kqyggq2V1H7wQj0/kJ3rMtfBBkfHeVhIeqjRJak8zrxmKF8FHSKUFNmx45F9n9kigyb
IkKmMXX27czmUE0NIGqqZq5kBxmH/dxp8H8mhqA9kWDE8Qul76BI28Ao9GcvE8vwnQLCq5kJauB6
+rcWkNnZac3sAy2PRDjZn7kjQbi8FawXhOvpageyNLnhFjmvLCvJnrMGqP9j1BOyLGOY6I8iOkV2
+igUKhqWKALH3qH3lppX86l/Z8IST0D+NLaDuPfcDCyik40olkLvk3z3h52eyGTkwlHjccYiOvZH
KXYGUU94rBFSiv8CPOuauc+JuhkwkPQ/D8+IchnHcTM7L/NKkoScdJwzpcSsGLidN6L1SegcbdNb
ciusdGaUPZyYrMItvtmW5Qkk+nMeZdxST6WScTN0WFqq7XgHwDma5Ltas4H6Pd2tkSNrWmVXBdTw
GaTsz0BGTKqma14Bh9iRr0ali+DCbqK2g19SxmmFvNp4uEXy2pgoBhaMvQv++bl28M15oBmlilnS
gs/OPnyeWKM1FcnTLy1cXXcUSOcFP73LrRCuwS11RmqoYa79JUIOaCLqsSYBjuRObXAb9rfpy4ue
1qPea05Cf2WLN8UWfcK/LryPYFz9tpfPbsHUo0GmxJ/aNm3EGFMazWNCqshE0iNWXUVzfCgN2/1m
R/AZQMuX40Wn90NscEwRUMhwOvoEwwNoQF6Ifq7HgX3nNlB/x+36K5py5aE/206a0Lt5xPUsRBrx
hcLp/NN+1CLrc9Yho1p86n2xjmIAhCZeZYDNsuIMisO9v70yVHkmvyPn3b4zvdhRz9dMdSbr1LZE
sAsmt4gq4n5ba5EkeUU9WHvqRgZboVbbiibiv1WlHZ8QTIEk+rGaoX/Ptv94tOWZAvH/kmtes1s0
VQijMNWhga2fMwuQqNBsq9nNafgdZAVrGDGruNwOZOYMKj5oulkE91Q8l6XOupuTrRzvEBGqHzGe
TVH3aFgA97Uhy2qXCPzuRVbm0fT89vGI27LGDyFb2InenjnAmH8eWv9wiREAz2ozFb1qo2+4ridW
KuBNaN1yCzzakgWUs4AXJH46W/yJBiUCt4fBQal0TZjhg5hkUINvvV5TcEMIg023Gf/dpI4+HoDJ
XHT4dRVgnQvd7oMWJ/lmlmAL2IesczcojIlNqkPfpPJSK3B7RmFigM0iFUIXpPFUHOgaH/OxE5ZF
DK2QDh6fCfm9CYgdPTXQ5urf/4D+bg1oKGEue/5FWHJRhFjo+ulTFiLar31WaCgutJcpgUAe/aYy
lwlLvSztITVkcS2mTEqnC351yNO2AS/35RTKcgvAVTyLSrjnP3/ULBOXVxT1h978Rt3jPOeWV/nl
4RvVHE7/M3n1hZHcaKGuIpZz4Q9r81chNj36aNnMzMAW4hAnMFNotbXfGB748PxJVF+8YUI5t3s2
9HM0J0mGoWgtLnjSkST6rYo3u58+P9Es6H+iQyEUa2pQze+/4pAkGcq1nJyuHdvpqP9N1ZRfFH44
lPATUW1d/2fHujQMkx4PL3lszhgS3I3Hzo5Z2PQCTDK+op17m18bzWIZviMlQabG1x300/F2maE9
+oTxKewYSY2JWaWghWx8vR/8n4VsIU4CW0Eyvnb0CcbfW9vIntvOn8XwmJ0txDhghnAOF6b24P7+
ogMhIHKRPOXVxJ1JDUf6z3zNZ5TgiIdKzciEt5AS7X/yx7cah4M+ONW4rdyaNnJaQZdDn7zD0HEo
2dZ1KeEMgEp8msL4d1FSK+BeWGWxaF/CbY2P75UtdJBqWxO8zgZz4ou0ZzzdZr3AQ8XLnoYKrB8z
zlpXvrms1ObsXUEccmiPBwwlwlpxgxoi92wMyEdbwWKE9IoLc+it1wBHyKwy+DnaQFXT6KkHIHy1
g/CgQKXfxfJ9e89o8SVrmgSSmEu7MdC2/8oHaQjqL7mR0sR9n8LV0vVuqf6isRof276qpoaOefqX
dGDh44lwTLT5/DKxBfWVT6CrlSSemz0EIPB5LMjt5+kD0ZWoBgRwQFaAuW05nDU8P7HnnadpUTNE
gSlb57I2fgAf6cBWiiLGJ/ZComRaDnoiiYO2xXIz6GIiIcvsFhmiwKEVJQ5nJ/euOPaKX1QWLzYu
fpZ6+f/1FlpxJv3B15PqvWafDUHbPCyttWPfi5kDEkGOe69YoQnyJ2/tIJga7E1cY1h8HRISUFHb
tvI19p8b/x+dLvS0CzFlhHZECe0DONraF8yEJp43FQDPjtnQW2vgBkpv0YRuNSdtq/00FjS+Z9FE
TKm61iBj+qx0zv++AMlRPx+xJBbsU+6I6MeKxp4Rjesxzv/Hr7CNhTChGXeodX/5K8XkRT2h+WnH
nnId2lVuZR8sEPN3hgUj4d/bl8kspztL9lXKPBgVVz8pUYMYWyXsEH6ebm7BxZtLc2eHUz2P+F2+
dKX37M19qOzFkBSVt5svV+aTWDHK23Bc6rC3h2M7Ie+6vZW8kuKcBF6KYg3ABpKngbmFHhhwZImg
vERtc2PGitgpw0HjqU34+skIppEIvPVKtzVljpGl5YArm/kAcGBK6+8sTh32g60EfM15Y0Lr4kfs
cbxoYDVen/Q/9l1k2hkNd21FN//RDztPcfVBBfknXbbCi90hcMOWXgPiIRVKmDmrpvsi1HWGLXUC
J2CA+31WL630k+E1gpohB8uD8gnAvrKj/KtlR/p7AiLfiARj4rKhkYZoUQpqafwwzdJzSxE3jGwt
ro7SV4C7CkIlFtiM4uA8g6YmrOgQfvi8umyI7BDgCIIc1ptdMReod/JNHOcJRePIf4xyiN+cUqg5
zevbE0qSj5XKpNIlRGmhhDahdcBHyk9WV0/Mq8E/t8/OEqwyBPSX+s3mqkDx79LuBHtKRVJjDu0P
pzO74eBDxWQJHx4eqMWGej+oamHfOAYIgIwyJZ5ptu2qI38ZNhiMOGbQtmlIH5M1TVqH9SuGwF23
pcRay9C4MspfwMY3YITuJJo7HpmzwQ7IRRDtvSqZaRAjskBSgByz/6N7NXQYoDyBxZ92KMbq56wn
0kft3HuXEW4ALEArQH6eONjhnPUMkjLMPT3r06J6l7Br/2vAYJJ4evoUSzSR+FcUPGwkfGCJ+iS6
2zJq9q/GxSxipobCM3GtMkt209+ol/CI6sTFYwz0bHTH2pI0Hd53f3GSqK2TANzLQqne6WZvnV+F
tF3qQIoGcGilIOL2Xb3gs+oW2lK8JqyexjCeJqZDcwm5IZ/4ED24K6/LT0PoR9YBTVU+wShIy4rL
lpqaKmrL4Pj0Eohycdw4xau4PTshxvEEYSnKzMkoOxHa1gtfvfRG343yUqgKOqy2bL8V/NZD1c/i
uHlw0aj2CNk55iyGCzGPzu+HheDyFT75e9DdTEZN3F4oUm92TLSUToUc9BCxWwJC8PmeM9tdQTc9
O4Z5Sr0jjw47igkRjwQ04c1Ri4S+91Btc9o3y8cm5wIdLhyZYtAU7QUX2BILBZNsN3fJzGIL3HEo
yDw7QcfEIY6P8MHJD/gSarskfkG/nEXX27uFKByPaW2vtsFGeHwZU7SN8ZzNQ0Qy/9CmaUHH7Tbo
FNukDiFyi4/sjvIdIMhfcnDEBiJFfaw8Yge+yU59PxjLZXVX1zy7MF14g+i3I53dPKIrEWw0oQ8+
NXZIpq1dcNorS2SmovtZbjRa6WwNKaqPvs7gC27UXmdIU50Zcc9z9Sq95gVfEwge0P8l/QupCrTT
tQv6/hGl2ZQLLrnHNqO7+24wiYjSQsIKVSD6UCjmv4qxPa57wlcfc+kRKiMtYbxiKH/g65BzN2sc
t0jlEnyOAenfmEp11ozLu6dLLz7vxk8Lx8ainmglMUQpyQfxFOj9LkDikJynrRm+0ZCebAZUeReP
loaUupp9JXHE/rYGPspXocVRPAirvjbtsFNPCLrOPCVIhVdOCLgSDi8fL0fJ1ZbuDGp8FVV1Gmq/
5CAqItFT/4tOd2sqY30RZyohv6V7KjVlWQ8GAsCCAYBtV5DpSqkMlqctiSt8wjmktIJyZVI0RF7I
+YNOZhX0F42eGue1NznZMUF0Ko1BWBZpPvlAEdip9Ap2r2NuXWhu1JSDcnvz1PIkOE6sH+N3E5cT
lGSoBqBFOafLdVskI7N7DQ5dAlbi2mMRO94xKPAPyB7Vsztsdd99kgUEKqgt6f5DFKUNsjVGi7C+
awHJfwdpqnE4Q14GJngSLeT0teOIjwlygRvvlnL887iO6opqlRxQMkp1sGYczq0NPj2+u04SCaIw
xtN6JjVWR2PbL9Is4B6De1hKwnuU8HUFKkbS6RL9PkzegYUz+IuxlSUVmMGZLEFLpITcU/5X1nUq
GS9E4F9qjmJFyQZy03RLQebiR1O9mmwueCTp3/fMQ8ZGXgmvGpGj76bzP40lZCaHbOh0KFEq0DNZ
LgXJ5keIbwwm+nPMXmYTd/0y1x19vHQeKcBy65eOAGqlyEgN16xyJY0Im8+FqlOuFofXG25I8HG1
ZjP1bRyB/tgPtjJehK75IbFxXkxCloziA9orJx77kDTMUyDe/qtm6u5JLsXT9AAMcNF4jcOj5Yb1
zGPsNexNSkHbnI3UuBAqJN+reRsonbeL7mJjJwugrMe+dFDitG5vXEUJIBlz73U1F1tiU1dMlJxZ
hZioRkdRk+xH7UfaY0NW3C+JhQ3MTq6DyN6qjL8ua9d3z6jkHjXOquOZXqqkQ5t0sB2Et1ttdslE
XiW492+BO5m6hW1acmF+Xcu+5lKzl84WOI/M35q3S5Jy1aoUowJZ85REhLS4+CXS+2WQJEdEGjBi
QVJuvyLaP7p3EBguwlQ7RavDkL7MWm10ovJNlKeMVOHSSqSMN0sSTcREWorqhJDXBrqICM05P9x4
UNx8TtNcSJfumf65S52mChAJIPDE4mOPc9L7ruvq9hFCJ6USbh5NF5Ahavsi1L26d/HPgh59chAU
/It6+3hRSC+o0mG4Dbj20UFiFKc7lERIodK9RDdGRwJaRTb40izGkSamWk/0Yd2SZAOLoH4YVnGa
DhxLlCxJUIPrec8uYBarqltCzonr+vQmaL0efXhTxo2Ivbmh0Ca2ybEwGI4Y3TgH14srF0CfXbfG
LGgUo1RBTKst/DvWbODSeNq+TZOjlwJA8gH+gr3Du8t4G+CE8jWyksMf6f+8C118zrfq6PjOPwXL
tLoKT6oBrI+s235Pt1kptiZDictn5DVC2FiUp2xXfVM6oP4Uc6NVlse9hZ8UtMPgGwSOGu+iaPZd
z+SznD1ep0K7ES8n/eanm4Jpf2f91ADcj4+wkt47yg4xV9BRw+KSSVFgBvdQwZyNxGQ2nwdGP/oq
PIwZI3QNI61F2b2LH+p/OEJCjjvGHZ7GGKXZRNyzBmHOofgCj/jCEPxRKrWCOIKwonYRw2j21Y7V
p8AEm8h5CjhhpRlPdM5N7h6bC1nTEvZ9IasWmQjnkJfwcaqBkgoPpovHFOP9fWTN/q5UllY1c3hV
bHBQEjifvy+gfTJs2h7olMjiZX7/sEsuq7bdEAsjeBhhStoAPqbP1LBBNIZWjpLbu9w9K3mbWT6e
xNOCRHe3TuvMow6OpOfXTLyqvgKrX1hd0btlkJu/Cg7jrFSBSY3WW0IeGeMqvJgmGkxVOAD8FLcE
YPl7pH4c9DUogycPznOxWCfLZdDY00e0bUyG1GpSVkhxXRA15nsOkteXPuPr4+nyEt/p9DLZkvzP
Wpel38UEYBCkRRqOW22n2Bovo5izv1p/9YBcYWaqN265qG3/QJOkrGuc/UoDeRmYrkeDkbziGhm+
6foRlGmxKPJClEjamK7OAUErNPJcmKNbKsLtYVQueAIJ48q83wsFM3mfl6bReXBheu68m2qETx7t
nfMAQKqh9rlBR/wDcuD5fALbM4a/sR7LfR1R98LMLx/JmWjG+73IZi13rI3NuywJRPFUuraWoCjn
lbjkEvxWG98eWEiSYlGLGBVBI9W+JCAYmq/iFKAJxmU657HcSJd3ONXQ5O3h73P6ysDBSIQ6AUyA
GycDZmlrPGm1Mfn3SJJtA1DftoWh8rmANnf5RPZW5CKcnRpV+4/bjMmgAgUcjnd13cRpGHL75HZv
YS7qaEoHmwmorMGC9vox5kxc5HleWtYdepnLa16aKEYqXBKiuV04AIwIJAT5U28mDMuVk2m1DgWL
53OLZESmU0jXcP3EEG2vz9GLtvyqYh+POBbBPJ5KbBjZF1GjH2vutHJtndoB2LmYdgx55xY+pMF2
w3gXlTd25Ny6nOomNtLa5nrCn1+O/BjcuV+SBMjys/fZkkkKUXbaV7sSjz7eFRquHPfIQIBX0blw
/2mWjunZdhHRcrRzxfbkw/e0hfRO/Oh1UIj15Z8ClpT6zVBXUFajxHr1t9iItfRBjFSzcPmjxnCh
9QX1gHgfekBK2z7WGGnGFTkXrOmyzMybxIRP65yxcpXqKWitZ9FZGyJuCpboeih0W9uoA+uoL/uo
pKk+wZsJtWDOjRcvQ6Hcn1geKhm8jULRSLm0zZpk8exsrcbWunbFXjGuUX+N2S46eq2pyHO4aI+r
wSEIjYc+SAtVnyl7iJrcDuoiw36Qo94jTJPK3KKyit8UIsEpPEc+Cp3G5TpQhnGM6kGUzuRnMj5x
IF5HusZvXNla3yUVpAuFHSoK1H2CrqKpMextCsxWUhIKR/KUfWqzPWVhiNlbwhwco4CN6gC+G2Mb
KdoVQM3gtFr3W+XGd0gzT0zBwt/AJXYL8WUpr2H9wRt+mCAEkvimAErcCtq8q68sTxmfBNUyzAZe
1B36Xc6p9TcHwm3EbE46y3nRowXme1n5PSxdFhDJwNkO6NYZ3k8Hqnhb23eSZS8teVeoTKoM8wUN
dl9CXvx5OQL4PL2SpS0uSrfcsS113bFCO7oqcS6xiHLosO3UPy9SxB8lyY83pmaoac7YZDLE+yyu
cvutxEfB/+ZNgdI0eJGEkCeXw/ab/4Oa8s61/mFNOgIt4kJ9ZCNzzWGTZGBTK7+pF+v9IaxXRNmp
LEsqQHj1TGw/Wv68YLCQoCf83aLzhYPcyVMTb8bvq2BWF/07SX1b0Y+iBVNsvCMlwGfboFoBe6mj
7onwY2wn7+veqsDE+N9BFeqJFjVw5Iazn+cSQUFGqW5VCN8Dpg0XbDeLycSurjJiyq/1pLKNSqKT
WOoCwrY6fvpS93ppFe+PWJNPtqo+fDpDG30BwTjjOaFAzEMxqE08OV+sJsZO3Ork5YxxNhjonHS3
bvjsydh0qzLfh2BtQJWtTfGe6Z9YnwhRDlUJA2sXxb9tz0+C5G2/unUC8LJATMBi27VA3sIJfJ1q
E6RpCt6mN2IHkAYSDcv2WjccvplkTS5GtKIgFFlYZ2mhxm87DfMpDGqZKCh25P1CZ04NQ/51d5Lg
9ovsYhiHGuYfYy8DQUt3/C53DAJbA9LrBdUoBBWxEZ3STkVA7TeVJyCrb2LzrI8j8jP81+f/y7ty
d0/HvMbw4iKsvtdRV7P1YY4LjDRV00ZfrYXJySdVtVd9N5pe6K07zIjw2vJtPICQIkp4zaQxgn7A
/ZByNWKjHfiGrcQ1ofMbSFP32xe3eQKV2bMzBX39f5jnjULD7jUOIuoVgJee/gd/WASI5aoXaEX5
gXbhu4YqM/6/D+fdhE7K2iPtxmprLOfViY3Psb1xvOSuju5x00i8wskYfprtONTjDykxSAWGtery
S4/45/kUcd7/BbtOt7wCgqy0jqXxJCQgkxKyKf3acrAR3xG3c6EeNcZ+5BCgiJl9RBkp4xhaNTaN
U9dPkK3uzGMUSf2CtUqEeG83urvjIQ==
`protect end_protected
